* NGSPICE file created from tt_um_essen.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_8 abstract view
.subckt sky130_fd_sc_hd__clkinv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_16 abstract view
.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

.subckt tt_um_essen VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4]
+ ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5]
+ uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5]
+ uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5]
+ uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7]
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1250/X m_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout554/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__and2b_2_B m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__a21o_2_A1/B1 sky130_fd_sc_hd__and2b_1
XFILLER_27_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout162_A fanout163/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_18_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout166/X m_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout619/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold22/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_50_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold491/A fanout57/X fanout69/X m_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__or2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout215_X fanout215/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__nor2_2_B fanout500/X hold1263/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B/A
+ hold616/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1 fanout450/X fanout456/X
+ fanout457/X fanout460/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1/X
+ sky130_fd_sc_hd__or4_1
XFILLER_50_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__xnor2_2_A hold1228/A hold599/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y
+ fanout39/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold351 hold351/A VGND VGND VPWR VPWR hold351/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold362 hold362/A VGND VGND VPWR VPWR hold362/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold340 hold340/A VGND VGND VPWR VPWR hold340/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout229/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout247/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhold395 hold395/A VGND VGND VPWR VPWR hold395/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold384 hold384/A VGND VGND VPWR VPWR hold384/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold373 hold373/A VGND VGND VPWR VPWR hold373/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_1430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout75_A fanout75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_5_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__a22o_2_A1 hold441/A fanout283/X
+ fanout406/X hold832/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1040 hold1040/A VGND VGND VPWR VPWR hold1040/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 hold1051/A VGND VGND VPWR VPWR hold1051/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 hold1062/A VGND VGND VPWR VPWR hold1062/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1084 hold1084/A VGND VGND VPWR VPWR hold1084/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold677/X m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold1073 hold1073/A VGND VGND VPWR VPWR hold1073/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1095 hold1095/A VGND VGND VPWR VPWR hold1095/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_16_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout30_X fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold39/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_70_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__or2_2_A_B fanout243/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold613/X hold654/X fanout562/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1270/A fanout44/X fanout72/X hold900/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1 m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold316/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout200/A m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout192/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_69_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_A1_N
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1256/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold124/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold831/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold576/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold1045/A fanout108/X fanout128/X hold407/A m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__or2_2_A_B fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XFILLER_75_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__a211oi_2_A1/Y m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2/Y
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X fanout406/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold228/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1135/X fanout228/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X_sky130_fd_sc_hd__xnor2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_A1 m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1086 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_A1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_S fanout155/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold512/X m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout297/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[13\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A hold659/X
+ VGND VGND VPWR VPWR hold658/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout157/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/D
+ fanout422/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_54_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout138 fanout139/X VGND VGND VPWR VPWR fanout138/X sky130_fd_sc_hd__clkbuf_4
Xfanout127 fanout127/A VGND VGND VPWR VPWR fanout127/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xfanout116 fanout119/A VGND VGND VPWR VPWR fanout116/X sky130_fd_sc_hd__buf_4
Xfanout105 fanout107/A VGND VGND VPWR VPWR fanout105/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold451/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A1_N
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout149 fanout151/X VGND VGND VPWR VPWR fanout149/X sky130_fd_sc_hd__buf_2
XANTENNA_m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1148/X fanout228/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout377_A fanout399/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.ll_q\[23\]_sky130_fd_sc_hd__or2_2_A hold371/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[23\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_43_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1122/A fanout92/X fanout148/X hold845/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X
+ hold185/A m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/B1 m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X/B1
+ fanout478/X ena_sky130_fd_sc_hd__or2_2_B/A VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[12\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold953/X VGND VGND VPWR VPWR hold1103/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__o22a_2_A2 fanout530/X hold368/A
+ m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__o22a_2_A2/B1 m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2
+ fanout288/X m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B/X fanout354/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold394/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1 hold403/A fanout278/X
+ fanout403/X hold655/A m_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__a22o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold332/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold314/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold170 hold170/A VGND VGND VPWR VPWR hold170/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_B
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/A
+ sky130_fd_sc_hd__nand2_1
Xhold192 hold192/A VGND VGND VPWR VPWR hold192/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 hold181/A VGND VGND VPWR VPWR hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/B
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/C m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ sky130_fd_sc_hd__a21bo_2
Xm_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_1 hold283/A m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout368/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout78_X fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__mux2_1_A0 hold311/X hold453/A
+ fanout605/X VGND VGND VPWR VPWR hold312/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_31_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold720/X fanout560/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout170/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold761/A sky130_fd_sc_hd__dfxtp_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_1 clkbuf_leaf_19_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1/D
+ VGND VGND VPWR VPWR uo_out[6] sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_leaf_46_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold293/X m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1/B1 m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout17/X hold162/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[6\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_15_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[12\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold926/X hold955/X fanout592/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X
+ hold1032/A fanout134/X m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X/A
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.g_buffer\[0\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_buffer\[21\].m_c_buf m_blake2.m_hash256.g_buffer\[21\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[21\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__o21ai_2_A1 hold1052/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout423/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_30_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout211/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or3b_2_B
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or3b_2_B/C_N
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or3b_2_B/X
+ sky130_fd_sc_hd__or3b_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_670 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[12\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1122/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold294/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/B1
+ sky130_fd_sc_hd__or2_1
XFILLER_29_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/B1
+ m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2/X
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_29_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_34_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_80_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[14\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1065/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_47_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_43_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1_A2
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
XANTENNA_fanout125_A fanout127/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__or2_2_B_A fanout486/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold112/X fanout317/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout494_A fanout500/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X
+ fanout107/X m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/B
+ sky130_fd_sc_hd__or4_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold546/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_58_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_X fanout282/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold599/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold946/A fanout84/X fanout140/X m_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_S fanout409/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[1\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold968/X hold626/X fanout560/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout260/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_67_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout38_A fanout39/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout86/X m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout107/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[10\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold671/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout214/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B fanout485/X hold212/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_23_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A hold349/A hold775/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold503/A fanout64/X fanout68/X hold758/A m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A0 hold81/A m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout534/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_1019 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[8\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold646/X m_blake2.m_hash256.m_matrix\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout588/X
+ VGND VGND VPWR VPWR hold647/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout278/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__mux2_1_A0 hold141/A m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout472/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout491 fanout493/X VGND VGND VPWR VPWR fanout491/X sky130_fd_sc_hd__buf_2
Xfanout480 fanout480/A VGND VGND VPWR VPWR fanout480/X sky130_fd_sc_hd__buf_4
XFILLER_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_Q
+ m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__or2_1
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__and2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ hold981/X VGND VGND VPWR VPWR hold980/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1 m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/C m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold928 hold928/A VGND VGND VPWR VPWR hold928/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold906 hold906/A VGND VGND VPWR VPWR hold906/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X
+ hold1097/A fanout91/X m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout393/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold140/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold917 hold917/A VGND VGND VPWR VPWR hold917/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_1_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload0/A sky130_fd_sc_hd__clkbuf_8
Xhold939 hold939/A VGND VGND VPWR VPWR hold939/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[9\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ hold1173/X VGND VGND VPWR VPWR hold1172/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold37/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_32_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__xor2_2_A hold870/A hold223/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold582/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__a22o_2_A1 hold1089/A fanout251/X
+ fanout170/X hold1185/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X/A2
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/B m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_buffer\[22\].m_y_buf m_blake2.m_hash256.g_buffer\[22\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[22\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__and2_2_B fanout439/X hold84/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold445/A fanout83/X fanout67/X m_blake2.m_hash256.m_matrix\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout110/X fanout134/X
+ hold1198/A m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout242_A fanout243/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__mux2_1_A0 hold97/A m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout508/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_io.m_config.ll_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold243/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout511/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout128_X fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2
+ fanout307/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A0 hold190/A m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout504/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout497_X fanout497/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/A3
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input2_X input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A
+ m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_matrix\[11\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold706/X hold732/X fanout586/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B fanout494/X hold111/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/A
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/B
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__nand3_2_B
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/B
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_matrix\[4\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold620/X m_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout575/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B_A fanout434/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold435/A fanout140/X fanout120/X hold720/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B fanout394/X fanout186/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/B1 sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.g_c_buf\[17\]_sky130_fd_sc_hd__a2111o_2_X m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout174/X m_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__o21a_2_A1/X
+ m_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__o21a_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[17\].m_c_buf/A sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_22_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_22_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_72_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout181/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold570/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X_X m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A0 hold41/A m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_20_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout64/X fanout36/X
+ hold890/A m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout200/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xhold703 hold703/A VGND VGND VPWR VPWR hold703/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[12\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1152/X m_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout551/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold714 hold714/A VGND VGND VPWR VPWR hold714/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold725 hold725/A VGND VGND VPWR VPWR hold725/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 hold736/A VGND VGND VPWR VPWR hold736/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 hold758/A VGND VGND VPWR VPWR hold758/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold747 hold747/A VGND VGND VPWR VPWR hold747/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold769 hold769/A VGND VGND VPWR VPWR hold769/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold656/A fanout146/X m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout107/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_44_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout192_A fanout192/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hash\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1 hash\[7\]_sky130_fd_sc_hd__and2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1 fanout462/X m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1/X sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__xnor2_2
XFILLER_26_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0 hold376/X m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold934/X hold980/A fanout545/X VGND VGND VPWR VPWR hold935/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout36/X fanout44/X
+ m_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1193/X hold988/X fanout590/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout412_X fanout412/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/X
+ m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__o21ai_2_A1/Y fanout268/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ fanout449/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__mux2_1_A1_S fanout323/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__xor2_2_B hold1265/A hold321/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1243/A fanout49/X fanout45/X hold727/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold63 hold63/A VGND VGND VPWR VPWR hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_5_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout60_X fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold74 hold74/A VGND VGND VPWR VPWR hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout343/X m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a21o_1
XFILLER_60_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_A_N_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31oi_2_Y/B1
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_3_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold96 hold96/A VGND VGND VPWR VPWR hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A VGND VGND VPWR VPWR hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[10\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold896/X hold744/X fanout567/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1198/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B fanout490/X hold152/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__xnor2_2_A hold342/A hold391/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1_B2 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__xnor2_2_B hold665/A hold506/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__mux2_1_A1 hold96/A m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout483/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2
+ fanout287/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1 hold532/A fanout381/X
+ fanout194/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A1
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A2
+ m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA_5 ANTENNA_5/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__xnor2_2_A hold922/A hold1174/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_50_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout260/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1_B1_N fanout409/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold36/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1120/A fanout50/X fanout74/X m_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__o2bb2a_2_A1_N m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout307/X fanout384/X hold348/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X
+ sky130_fd_sc_hd__o2bb2a_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A fanout449/A fanout458/X
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/C VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold100/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold511 hold511/A VGND VGND VPWR VPWR hold511/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold500 hold500/A VGND VGND VPWR VPWR hold500/X sky130_fd_sc_hd__dlygate4sd3_1
Xhash\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hash\[6\]_sky130_fd_sc_hd__or2_2_B/B fanout335/X VGND VGND VPWR VPWR hash\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold522 hold522/A VGND VGND VPWR VPWR hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout205_A fanout208/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold533 hold533/A VGND VGND VPWR VPWR hold533/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[15\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold886/X hold300/X fanout574/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold544 hold544/A VGND VGND VPWR VPWR hold544/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 hold577/A VGND VGND VPWR VPWR hold577/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold555 hold555/A VGND VGND VPWR VPWR hold555/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ sky130_fd_sc_hd__and2b_1
Xhold566 hold566/A VGND VGND VPWR VPWR hold566/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold588 hold588/A VGND VGND VPWR VPWR hold588/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B_A fanout492/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold599 hold599/A VGND VGND VPWR VPWR hold599/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout286/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o22a_1
Xhold1200 hold1200/A VGND VGND VPWR VPWR hold1200/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout195_X fanout195/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1222 hold1222/A VGND VGND VPWR VPWR hold1222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1211 hold1211/A VGND VGND VPWR VPWR hold1211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1233 hold1233/A VGND VGND VPWR VPWR hold1233/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1255 hold1255/A VGND VGND VPWR VPWR hold1255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1244 hold1244/A VGND VGND VPWR VPWR hold1244/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__xnor2_2_A hold284/A hold1244/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold1266 hold1266/A VGND VGND VPWR VPWR hold1266/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold833/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_2_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold356/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__or2_2_A hold204/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold511/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A0 hold174/A m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout508/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_B2
+ fanout267/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_A1
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout285/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_8_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XFILLER_76_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A_A m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X
+ hold444/A fanout345/X fanout181/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold261/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1247/X m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout153/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X/A1
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D/Y
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/A
+ sky130_fd_sc_hd__a21bo_2
XFILLER_60_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout18/X m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[9\].m_y_buf/A sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold71/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__a22o_2_A1 hold715/A fanout292/X
+ fanout287/X hold616/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ hold310/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1/X
+ sky130_fd_sc_hd__o311a_1
Xfanout309 fanout314/X VGND VGND VPWR VPWR fanout309/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold704/X m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout294/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A0 hold151/A m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout516/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout233/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold573/X fanout162/X m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/A
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/C
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/X
+ sky130_fd_sc_hd__or4_1
XFILLER_54_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__a22o_2_A1_A1 m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_18_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__a22o_2_A1 hold337/A fanout192/X
+ fanout200/X hold488/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout155_A fanout156/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout322_A fanout323/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1198/X hold1057/X fanout586/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout110_X fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__a22o_2_A1 hold432/A fanout187/X
+ fanout195/X hold860/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout269/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout208_X fanout208/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/B1
+ sky130_fd_sc_hd__nand2b_1
Xm_blake2.m_hash256.m_matrix\[10\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[10\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1076/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ fanout614/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xhold352 hold352/A VGND VGND VPWR VPWR hold352/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[0\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/B2 hold893/A fanout558/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold341 hold341/A VGND VGND VPWR VPWR hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 hold330/A VGND VGND VPWR VPWR hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 hold396/A VGND VGND VPWR VPWR hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 hold385/A VGND VGND VPWR VPWR hold385/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 hold374/A VGND VGND VPWR VPWR hold374/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout289/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold363 hold363/A VGND VGND VPWR VPWR hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout203/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout68_A fanout71/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1030 hold1030/A VGND VGND VPWR VPWR hold1030/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__o21a_2
Xhold1041 hold1041/A VGND VGND VPWR VPWR hold1041/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1052 hold1052/A VGND VGND VPWR VPWR hold1052/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 hold1074/A VGND VGND VPWR VPWR hold1074/X sky130_fd_sc_hd__dlygate4sd3_1
Xdata\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X data\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1047/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1085 hold1085/A VGND VGND VPWR VPWR hold1085/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1063 hold1063/A VGND VGND VPWR VPWR hold1063/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1096 hold1096/A VGND VGND VPWR VPWR hold1096/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A_B fanout487/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_900 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xdata\[6\]_sky130_fd_sc_hd__mux2_1_A1 data\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold199/X
+ fanout579/X VGND VGND VPWR VPWR data\[6\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A1
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A2
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A3
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/B sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.m_matrix\[7\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold998/X m_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout587/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_clkbuf_leaf_5_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1166/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout200/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2
+ fanout274/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold70/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__or2_2_A/A fanout161/X m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout614/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_68_1364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold885/A fanout140/X fanout92/X m_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhash\[0\]_sky130_fd_sc_hd__or2_2_B fanout483/X hash\[0\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR hash\[0\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__and2_1
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[13\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.v_q\[13\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold915/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A_A
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1207/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold260/X m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_1302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/A1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ sky130_fd_sc_hd__a21boi_4
XFILLER_33_900 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__a21oi_2_A1 hold282/A fanout282/X
+ m_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__a22o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__a21oi_2_A1/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1 m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1/A2
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_33_988 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_45_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1092 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1019/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold838/X m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout418/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_B1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__nor3_2_Y
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__nor3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/D m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xfanout106 fanout107/A VGND VGND VPWR VPWR fanout106/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout417/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout117 fanout119/A VGND VGND VPWR VPWR fanout117/X sky130_fd_sc_hd__buf_2
Xfanout128 fanout131/A VGND VGND VPWR VPWR fanout128/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xfanout139 fanout139/A VGND VGND VPWR VPWR fanout139/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout18/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout272_A fanout273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X
+ fanout192/X m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o2bb2a_1
Xm_blake2.m_hash256.m_matrix\[11\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold654/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout537_A fanout538/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_X fanout158/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold467/X m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_A
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout190/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold485/X m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout297/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold459/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout412/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold160 hold160/A VGND VGND VPWR VPWR hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 hold171/A VGND VGND VPWR VPWR hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_C
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold193 hold193/A VGND VGND VPWR VPWR hold193/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[3\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold491/X hold400/X fanout572/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold182 hold182/A VGND VGND VPWR VPWR hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold78/A m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout530/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[12\]\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold965/X fanout227/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[0\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ hold684/X VGND VGND VPWR VPWR hold683/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout176/A fanout273/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
XFILLER_74_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/A2
+ sky130_fd_sc_hd__and3b_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_2 clkbuf_leaf_19_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2/D
+ VGND VGND VPWR VPWR uo_out[5] sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__a21o_2_A1_A2 fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_2
XFILLER_27_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_42_730 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[15\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ data\[0\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold275/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[3\]_sky130_fd_sc_hd__mux2_1_A1_S fanout228/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold60/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_S fanout222/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout155/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold322/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ hold544/X VGND VGND VPWR VPWR hold543/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_buffer\[25\].m_c_buf m_blake2.m_hash256.g_buffer\[25\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[25\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout168/X m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout621/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1 hold829/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout427/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_10_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold525/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold400/A fanout133/X fanout121/X hold300/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_1058 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B/X sky130_fd_sc_hd__and2b_1
XFILLER_49_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout41/X fanout37/X
+ hold1080/A m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_34_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold798/A fanout38/X fanout46/X m_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout186/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_37_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[29\]_sky130_fd_sc_hd__o21a_2_A1 hold448/A fanout386/X
+ fanout170/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.m_matrix\[4\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1078/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[8\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[8\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold726/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[11\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1175/X hold1231/A fanout552/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or3_2_A_1 fanout450/X fanout456/X
+ fanout462/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/D
+ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_47_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__a21o_2_A1 hold273/X fanout321/X
+ m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_43_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[8\]\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold793/X fanout222/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_43_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout118_A fanout119/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1084/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__a22oi_2_B2_B2 m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A fanout489/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2_B1_sky130_fd_sc_hd__nand2_2_Y_A
+ fanout463/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_60_1456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout275_X fanout275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_X fanout442/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a31o_2_A2
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.m_matrix\[8\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[8\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold950/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o32a_2_X
+ fanout498/X m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A/Y fanout274/X
+ m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o32a_1
XANTENNA_clkbuf_3_5_0_clk_X clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold211/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold157/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold81/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout90_X fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold141/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_S fanout302/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout476/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout492 fanout493/X VGND VGND VPWR VPWR fanout492/X sky130_fd_sc_hd__buf_2
Xfanout481 fanout482/X VGND VGND VPWR VPWR fanout481/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout470 fanout471/X VGND VGND VPWR VPWR fanout470/X sky130_fd_sc_hd__dlymetal6s2s_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_B1_sky130_fd_sc_hd__or3b_2_X
+ fanout458/X fanout460/X fanout468/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X/B1
+ sky130_fd_sc_hd__or3b_1
XFILLER_24_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout280/X m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout287/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A hold374/A m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_30_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o21ai_1
Xhold907 hold907/A VGND VGND VPWR VPWR hold907/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_A_N_B
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold918 hold918/A VGND VGND VPWR VPWR hold918/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold929 hold929/A VGND VGND VPWR VPWR hold929/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__or4_2_B_D_sky130_fd_sc_hd__or4_2_X
+ hold1/A hold5/A hold2/A fanout308/X VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__or4_2_B/D
+ sky130_fd_sc_hd__or4_1
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A hold310/A m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1 hold271/A m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout375/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_36_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X/B
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_9_1036 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/A
+ sky130_fd_sc_hd__inv_2
XFILLER_56_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout551/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold123/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[10\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1167/X hold1187/A fanout594/X VGND VGND VPWR VPWR hold1168/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold939/X fanout557/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X
+ fanout111/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[26\].m_y_buf m_blake2.m_hash256.g_buffer\[26\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[26\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold188/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout235_A fanout236/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A2
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/A2
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout402_A fanout403/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__a21o_2_A1 hold45/X fanout327/X
+ m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__o21ba_2_X
+ m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y/A m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__o21ba_1
Xm_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_45_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout414/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__o22a_2_A2/B1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold190/X fanout309/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__a31o_2_A3 fanout472/X fanout476/X
+ hold518/A fanout366/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout347/X m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X fanout256/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout130/X
+ fanout118/X hold1117/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_67_clk clkload0/A VGND VGND VPWR VPWR clkload11/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.g_buffer\[5\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout50_A fanout51/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout520/X m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_891 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold359/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__mux2_1_A0 hold10/A m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout526/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_76_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout186/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__xnor2_2_A hold314/A hold951/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__and2_2_B fanout428/X hold210/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_30_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__a221o_2_B2_C1 fanout268/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_clk clkload3/A VGND VGND VPWR VPWR clkbuf_leaf_58_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
XFILLER_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout258/X m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout394/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold177/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__xnor2_2_A_B m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3
+ fanout470/X fanout475/X m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout346/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold41/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold737 hold737/A VGND VGND VPWR VPWR hold737/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 hold726/A VGND VGND VPWR VPWR hold726/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold704 hold704/A VGND VGND VPWR VPWR hold704/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 hold715/A VGND VGND VPWR VPWR hold715/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ hold1261/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 fanout240/X hold268/A
+ m_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XANTENNA_m_blake2.m_hash256.m_matrix\[3\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold748 hold748/A VGND VGND VPWR VPWR hold748/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold959/A fanout116/X fanout148/X m_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout417/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold759 hold759/A VGND VGND VPWR VPWR hold759/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__o2bb2a_2_A1_N_A2_N fanout307/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout185_A fanout186/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_49_clk clkload2/A VGND VGND VPWR VPWR clkload20/A sky130_fd_sc_hd__clkbuf_8
Xm_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__o22a_2_A1_A2 m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1/Y m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__a21oi_2_B1 m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold216/A VGND VGND VPWR VPWR m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_68_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.g_buffer\[11\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__a211o_2_A1 hold506/A fanout279/X
+ m_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__a22o_2_A1/X fanout372/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold730/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout617_A fanout621/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout140_X fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X fanout445/X m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A0 hold274/A m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout501/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout222/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/A
+ hold468/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B fanout426/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y
+ m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1150/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout98_A fanout99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_1_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A VGND VGND VPWR VPWR hold64/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout256/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__xnor2_2_A hold350/A hold1135/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1033/X fanout555/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold97 hold97/A VGND VGND VPWR VPWR hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A VGND VGND VPWR VPWR hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xhold75 hold75/A VGND VGND VPWR VPWR hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout50/X fanout46/X
+ hold849/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1_A2 m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_0_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_3_0_0_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
XFILLER_40_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1
+ fanout286/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2_sky130_fd_sc_hd__nor2_2_Y_A
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_74_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__or2_2_B_A fanout478/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 ANTENNA_6/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/D
+ m_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout229/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__xnor2_2_A hold1087/A hold464/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout25/X fanout29/X
+ m_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__a21oi_2_B1_B1 m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nand2b_2_Y_B
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_6_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or2_2_B fanout456/X hold1180/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/C sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_50_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A0 hold60/A m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/A2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ hold1160/X m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout425/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2
+ fanout266/X m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__nand2_2_B/Y
+ fanout400/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ sky130_fd_sc_hd__o22ai_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload23/A m_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_76_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y
+ hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__xnor2_2_B hold598/A hold479/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold501 hold501/A VGND VGND VPWR VPWR hold501/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 hold534/A VGND VGND VPWR VPWR hold534/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold523 hold523/A VGND VGND VPWR VPWR hold523/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold512 hold512/A VGND VGND VPWR VPWR hold512/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout100_A fanout103/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold545 hold545/A VGND VGND VPWR VPWR hold545/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/C
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__o21ai_2
Xhold578 hold578/A VGND VGND VPWR VPWR hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold567 hold567/A VGND VGND VPWR VPWR hold567/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 hold556/A VGND VGND VPWR VPWR hold556/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__and3_2_B_B
+ m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold589 hold589/A VGND VGND VPWR VPWR hold589/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B_B m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold295/A m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__or2_2_B/X fanout382/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1234 hold1234/A VGND VGND VPWR VPWR hold1234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1212 hold1212/A VGND VGND VPWR VPWR hold1212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1201 hold1201/A VGND VGND VPWR VPWR hold1201/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1223 hold1223/A VGND VGND VPWR VPWR hold1223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1256 hold1256/A VGND VGND VPWR VPWR hold1256/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1245 hold1245/A VGND VGND VPWR VPWR hold1245/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout188_X fanout188/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1267 hold1267/A VGND VGND VPWR VPWR hold1267/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout62/X fanout30/X
+ m_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1164/A fanout62/X fanout38/X hold1222/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout355_X fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1061/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout258/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_26_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout303/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold966/X fanout221/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold174/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold727/X hold1178/A fanout576/X VGND VGND VPWR VPWR hold728/A sky130_fd_sc_hd__mux2_1
XFILLER_16_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X
+ m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_S fanout153/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_S fanout158/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N/X
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__a31o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1 m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout426/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout351/X m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X fanout258/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1067/X fanout593/X
+ VGND VGND VPWR VPWR hold1068/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[5\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__a32o_2_A1_A3 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B fanout429/X hold222/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_64_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold777/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[9\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold880/X hold817/X fanout544/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold890/X hold768/A fanout553/X VGND VGND VPWR VPWR hold891/A sky130_fd_sc_hd__mux2_1
XFILLER_17_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__xor2_2_A hold488/A hold1055/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1241/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold439/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold914/X fanout592/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__or2_2_A hold643/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__o21a_2_A1 hold966/A fanout366/X
+ fanout254/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_1 hold254/A m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout374/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold629/X m_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout551/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__and3_2_A hold306/A fanout465/X fanout376/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X
+ fanout106/X m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X/B
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A/B
+ sky130_fd_sc_hd__or3_2
XTAP_TAPCELL_ROW_52_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X_A2 fanout174/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold192/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_52_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__inv_2_A fanout474/X VGND VGND VPWR
+ VPWR fanout408/A sky130_fd_sc_hd__inv_2
XFILLER_41_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1110/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold151/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/X fanout609/X input8/X VGND VGND VPWR VPWR m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
XFILLER_35_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_62_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_23_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_18_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout360/X m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ fanout179/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__and3b_2_X
+ fanout468/X fanout469/X fanout474/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ sky130_fd_sc_hd__and3b_2
XANTENNA_fanout148_A fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[6\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[12\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold636/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__a22o_2_A1 hold618/A fanout295/X
+ fanout283/X hold666/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xhold320 hold320/A VGND VGND VPWR VPWR hold320/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold342 hold342/A VGND VGND VPWR VPWR hold342/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold714/X fanout226/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout103_X fanout103/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1179/A sky130_fd_sc_hd__dfxtp_1
Xhold331 hold331/A VGND VGND VPWR VPWR hold331/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold353 hold353/A VGND VGND VPWR VPWR hold353/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
Xhold364 hold364/A VGND VGND VPWR VPWR hold364/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 hold386/A VGND VGND VPWR VPWR hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 hold375/A VGND VGND VPWR VPWR hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 hold397/A VGND VGND VPWR VPWR hold397/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
XFILLER_24_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1042 hold1042/A VGND VGND VPWR VPWR hold1042/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 hold1031/A VGND VGND VPWR VPWR hold1031/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout472_X fanout472/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1020 hold1020/A VGND VGND VPWR VPWR hold1020/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__mux2_1_A0 hold76/A m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold389/A sky130_fd_sc_hd__dfxtp_1
Xhold1064 hold1064/A VGND VGND VPWR VPWR hold1064/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1075 hold1075/A VGND VGND VPWR VPWR hold1075/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__a211oi_2_A1_A2 fanout288/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1053 hold1053/A VGND VGND VPWR VPWR hold1053/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[10\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold665/X m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout234/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold1097 hold1097/A VGND VGND VPWR VPWR hold1097/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 hold1086/A VGND VGND VPWR VPWR hold1086/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold1016/A fanout85/X fanout133/X hold1000/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/B
+ m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout415/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout16_X fanout16/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3
+ fanout451/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C/X
+ fanout444/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3/X
+ sky130_fd_sc_hd__o31a_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout91/X
+ fanout135/X hold954/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/B2
+ hold909/X fanout577/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__a22o_2_A1 hold374/A fanout191/X
+ fanout199/X hold788/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_B_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/D
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/B
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold272/X m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout232/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_S fanout412/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold464/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout358/X m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__a22o_2_A1/X fanout179/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout55/X
+ fanout82/X m_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.g_buffer\[5\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_51_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold519/X m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[12\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold424/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1046/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold420/A m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout380/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__xor2_2_A hold799/A hold942/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_41_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_41_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold318/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold979/X fanout219/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/Y m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_Y
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A0 hold42/A m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout508/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold592/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[14\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A hold531/X
+ VGND VGND VPWR VPWR hold530/A sky130_fd_sc_hd__dfxtp_1
Xfanout107 fanout107/A VGND VGND VPWR VPWR fanout107/X sky130_fd_sc_hd__clkbuf_2
Xfanout118 fanout119/A VGND VGND VPWR VPWR fanout118/X sky130_fd_sc_hd__clkbuf_4
Xfanout129 fanout131/A VGND VGND VPWR VPWR fanout129/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1199/X
+ fanout558/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1
+ fanout285/X m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout279/X fanout350/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_68_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold612/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout299/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1
+ fanout286/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold507/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A/B fanout206/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold796/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout432_A fanout434/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold927/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/X m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold1214/X fanout218/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[20\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XANTENNA_fanout220_X fanout220/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold753/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_30_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold836/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold546/X m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1015/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold207/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1147/A fanout126/X fanout90/X hold1130/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xhold150 hold150/A VGND VGND VPWR VPWR hold150/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__a221o_2_A1 hold1142/A m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ m_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__or2_2_A/X fanout171/X m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__o21a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[10\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a221o_1
Xhold161 hold161/A VGND VGND VPWR VPWR hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_2
Xhold194 hold194/A VGND VGND VPWR VPWR hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A VGND VGND VPWR VPWR hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold172 hold172/A VGND VGND VPWR VPWR hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold78/X fanout335/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold888/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout80_A fanout83/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold748/A fanout117/X fanout149/X hold421/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold428/X m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__a221o_2_A1 hold1225/A fanout352/X
+ fanout264/X m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout393/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_1_0_clk_X clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__nor2_2_B fanout488/X hold250/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__a21bo_2_A2
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__a21bo_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_3 clkbuf_leaf_20_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3/D
+ VGND VGND VPWR VPWR uo_out[4] sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[5\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold794/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_33_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold904/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__xnor2_2_A hold619/A hold730/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XFILLER_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.g_buffer\[13\].m_c_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__mux2_1_A0 hold169/A m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout523/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold986/X fanout164/X m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_matrix\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold693/X hold553/X fanout556/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[11\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[11\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1040/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__mux2_1_A0 hold93/A m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold189/X m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout299/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_A_N
+ m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout170/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout251/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[29\].m_c_buf m_blake2.m_hash256.g_buffer\[29\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[29\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold998/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__nand2b_2
Xm_blake2.m_hash256.m_matrix\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1111/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ fanout461/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/X fanout612/X VGND VGND VPWR VPWR
+ m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_34_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout291/X m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_64_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[15\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ data\[6\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR data\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold88/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[9\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[9\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1213/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_43_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B/A
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B/Y
+ sky130_fd_sc_hd__nor3_1
XFILLER_53_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold418/X m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout156/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[28\]_sky130_fd_sc_hd__or2_2_A hold1064/A fanout247/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[28\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B fanout490/X hold89/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout382_A fanout385/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold233/X fanout165/X m_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout268_X fanout268/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2
+ fanout168/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_X fanout170/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold871/A fanout28/X m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/B2 hold1224/A m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout435_X fanout435/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ m_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout612/X VGND VGND VPWR VPWR m_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A0 hold39/A m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1183/X hold1248/A fanout580/X VGND VGND VPWR VPWR hold1184/A sky130_fd_sc_hd__mux2_1
XFILLER_30_1272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_2_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout35/X fanout47/X
+ hold725/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X
+ hold1264/A fanout27/X m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout23/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold704/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xfanout493 fanout494/X VGND VGND VPWR VPWR fanout493/X sky130_fd_sc_hd__clkbuf_2
Xfanout482 hold1075/A VGND VGND VPWR VPWR fanout482/X sky130_fd_sc_hd__buf_2
Xfanout460 fanout460/A VGND VGND VPWR VPWR fanout460/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout471 fanout472/X VGND VGND VPWR VPWR fanout471/X sky130_fd_sc_hd__buf_4
XFILLER_4_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X_A2 fanout275/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and2_2_A/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[8\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold407/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__a221o_2_A1 hold806/A fanout275/X
+ fanout176/X m_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__or2_2_A/X fanout271/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold908 hold908/A VGND VGND VPWR VPWR hold908/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__a21oi_1
Xhold919 hold919/A VGND VGND VPWR VPWR hold919/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_36_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_A1
+ fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1048 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout295/X m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B/X m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout406/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold928/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_65_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout422/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_53_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_S
+ fanout435/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout201/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout130_A fanout131/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_A fanout228/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A_Y m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1 fanout454/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1/X sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2
+ fanout257/X m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ fanout397/X fanout179/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0 hold1055/X m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ hold535/X fanout276/X m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout415/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold424/A fanout82/X fanout66/X m_blake2.m_hash256.m_matrix\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__a22o_2_B2 hold1161/A fanout259/X fanout304/X
+ hold605/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout385_X fanout385/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__or2_2_B fanout497/X hold188/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_25_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1242/X fanout566/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold139/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1 m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/B2
+ fanout100/X m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/Y sky130_fd_sc_hd__o22ai_4
Xm_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_A
+ fanout408/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1/X m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_22_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout422/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1136/X fanout544/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__mux2_1_A1_S fanout330/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__a31o_2_B1 hold1260/A
+ m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B
+ m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
Xm_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout290 fanout291/X VGND VGND VPWR VPWR fanout290/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__xnor2_2_A hold293/A hold851/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_47_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_76_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__xor2_2_A hold805/A hold247/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/A2
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/B1
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout192/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__xnor2_2_A hold525/A hold603/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold705 hold705/A VGND VGND VPWR VPWR hold705/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold582/A fanout114/X m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A2
+ sky130_fd_sc_hd__a2111o_1
Xhold727 hold727/A VGND VGND VPWR VPWR hold727/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 hold716/A VGND VGND VPWR VPWR hold716/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__or2_2_A hold201/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xhold738 hold738/A VGND VGND VPWR VPWR hold738/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold749 hold749/A VGND VGND VPWR VPWR hold749/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__o211a_2_A1_A1 m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A1_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_X clkload14/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold651/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout178_A fanout180/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold344/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__nor2_4
XFILLER_0_1354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout345_A fanout346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold122/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout273/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold274/X fanout309/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1111/A fanout51/X fanout46/X hold718/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_io.m_block_data.data_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ hold6/A m_io.data_v_early_sky130_fd_sc_hd__and3_2_C/X m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout300_X fanout300/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__or2_2_B fanout486/X hold864/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1058/X hold1130/A fanout583/X VGND VGND VPWR VPWR hold1059/A sky130_fd_sc_hd__mux2_1
XFILLER_62_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xor2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold65 hold65/A VGND VGND VPWR VPWR hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold87 hold87/A VGND VGND VPWR VPWR hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A VGND VGND VPWR VPWR hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[7\]_sky130_fd_sc_hd__or2_2_A hold1092/A fanout393/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[7\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhold98 hold98/A VGND VGND VPWR VPWR hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout551/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A0 hold386/A m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout46_X fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__and2_2_B fanout429/X hold1012/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N/Y
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1/Y
+ sky130_fd_sc_hd__a21boi_1
XFILLER_73_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2_sky130_fd_sc_hd__nor2_2_Y_B
+ m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_X m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2 m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/A1
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/A2 m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/A3
+ fanout102/X hold311/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/X
+ sky130_fd_sc_hd__o32a_2
XANTENNA_7 ANTENNA_8/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_4_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout413/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__nand2_1
XFILLER_80_1449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold115/A sky130_fd_sc_hd__dfxtp_1
XFILLER_39_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_50_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold60/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B/A
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_1/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B/Y
+ sky130_fd_sc_hd__nor4_1
Xm_blake2.m_hash256.m_matrix\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1101/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B/X m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_clkbuf_leaf_44_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XFILLER_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__nand2b_2_B fanout466/X fanout462/X
+ VGND VGND VPWR VPWR fanout361/A sky130_fd_sc_hd__nand2b_4
XFILLER_31_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__xnor2_1
XFILLER_31_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1227/X
+ fanout558/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/B1
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_11_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_59_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout448/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xhold502 hold502/A VGND VGND VPWR VPWR hold502/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A hold406/A m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
Xhold535 hold535/A VGND VGND VPWR VPWR hold535/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold524 hold524/A VGND VGND VPWR VPWR hold524/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 hold513/A VGND VGND VPWR VPWR hold513/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 hold546/A VGND VGND VPWR VPWR hold546/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 hold568/A VGND VGND VPWR VPWR hold568/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold557 hold557/A VGND VGND VPWR VPWR hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 hold579/A VGND VGND VPWR VPWR hold579/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_58_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout295_A fanout295/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1213 hold1213/A VGND VGND VPWR VPWR hold1213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1224 hold1224/A VGND VGND VPWR VPWR hold1224/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/A
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ sky130_fd_sc_hd__or3_1
Xhold1202 hold1202/A VGND VGND VPWR VPWR hold1202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1246 hold1246/A VGND VGND VPWR VPWR hold1246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1235 hold1235/A VGND VGND VPWR VPWR hold1235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1257 hold255/A VGND VGND VPWR VPWR hold1257/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1268 hold216/A VGND VGND VPWR VPWR hold1268/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_A fanout615/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout250_X fanout250/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_A
+ fanout269/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_24_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout17/X hold1233/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[23\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_S fanout420/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_700 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout291/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__nand2_2_B/Y
+ fanout400/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ sky130_fd_sc_hd__o22ai_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_B1
+ fanout103/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout18/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B_A fanout489/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1026/A fanout56/X fanout72/X hold1078/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold974/A fanout115/X fanout146/X m_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2/A1
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__nor2_2_B fanout491/X hold173/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_60_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/B1
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X/A sky130_fd_sc_hd__nand2b_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X/A2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X/B1
+ hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_73_1242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0_S fanout299/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A fanout472/X fanout476/X
+ VGND VGND VPWR VPWR fanout406/A sky130_fd_sc_hd__nor2_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_B2 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold556/X m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout116/X
+ fanout144/X hold456/A m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/B
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A
+ hold843/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[4\]_sky130_fd_sc_hd__mux2_1_A1_S fanout228/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_S fanout224/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__o41a_2_X
+ fanout455/X fanout459/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D/C
+ sky130_fd_sc_hd__o41a_1
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout67/X
+ fanout79/X hold790/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold327/X m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout316/X VGND VGND VPWR VPWR hash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold455/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout210_A fanout211/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ hold1217/X m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/A_N
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__o311a_2_A1/X VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xhold310 hold310/A VGND VGND VPWR VPWR hold310/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout295/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_S fanout231/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold343 hold343/A VGND VGND VPWR VPWR hold343/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 hold332/A VGND VGND VPWR VPWR hold332/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold321/A VGND VGND VPWR VPWR hold321/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2
+ fanout406/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Left_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold832/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout241/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhold376 hold376/A VGND VGND VPWR VPWR hold376/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 hold387/A VGND VGND VPWR VPWR hold387/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold354 hold354/A VGND VGND VPWR VPWR hold354/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 hold365/A VGND VGND VPWR VPWR hold365/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xhold398 hold398/A VGND VGND VPWR VPWR hold398/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold273/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[10\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[10\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold1137/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold446/X m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold1032 hold1032/A VGND VGND VPWR VPWR hold1032/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1010 hold1010/A VGND VGND VPWR VPWR hold1010/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1021 hold1021/A VGND VGND VPWR VPWR hold1021/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1054 hold1054/A VGND VGND VPWR VPWR hold1054/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 hold1043/A VGND VGND VPWR VPWR hold1043/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout465_X fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1076 hold1076/A VGND VGND VPWR VPWR hold1076/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_39_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A/B
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
Xhold1065 hold1065/A VGND VGND VPWR VPWR hold1065/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1098 hold1098/A VGND VGND VPWR VPWR hold1098/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1087 hold1087/A VGND VGND VPWR VPWR hold1087/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold441/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1094/X hold1115/A fanout554/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A hold186/X
+ VGND VGND VPWR VPWR hold216/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold1174/X m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[13\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1250/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ hold163/X VGND VGND VPWR VPWR hold162/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold858/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold370/A m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__or2_2_B/X fanout381/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XFILLER_10_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[0\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1004/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout192/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[23\]_sky130_fd_sc_hd__o311a_2_X fanout477/X hold1230/A
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.g_c_buf\[23\]_sky130_fd_sc_hd__o311a_2_X/B1
+ fanout355/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[23\].m_c_buf/A sky130_fd_sc_hd__o311a_1
XFILLER_68_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[12\]\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1163/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold295/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_69_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/B fanout370/X fanout185/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X/B1 sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__and4_2_C m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1245/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/D
+ sky130_fd_sc_hd__and4_2
Xm_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__a22o_2_A1 hold628/A fanout169/X
+ fanout171/X hold1214/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[2\]_sky130_fd_sc_hd__a211o_2_X/A2
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[15\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ data\[5\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR data\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold940/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold598/X m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold905/X m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout156/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold568/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[2\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ hold850/X VGND VGND VPWR VPWR hold849/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold373/X m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout414/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a311oi_2_Y
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/A m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X/B
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2/X
+ VGND VGND VPWR VPWR ANTENNA_6/DIODE sky130_fd_sc_hd__a311oi_4
XFILLER_73_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold313/X fanout216/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold420/X fanout216/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold164/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B_A fanout485/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ hold422/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold42/X fanout317/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout607/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout301/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout119 fanout119/A VGND VGND VPWR VPWR fanout119/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold256/X m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout232/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold625/X VGND VGND VPWR VPWR hold624/A sky130_fd_sc_hd__dfxtp_1
Xfanout108 fanout111/A VGND VGND VPWR VPWR fanout108/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[8\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1203/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold667/A fanout53/X m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__a21o_2_A1 hold17/X fanout339/X
+ m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y
+ fanout186/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout221/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1238/X hold1209/X fanout584/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout221/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold781/A fanout50/X fanout74/X hold1193/A m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X_B1 m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A fanout258/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout160_A fanout160/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[12\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1227/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1003/X hold937/X fanout557/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout425_A fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold298/A m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout383/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout418/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ hold723/X VGND VGND VPWR VPWR hold722/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout124/X
+ fanout120/X data\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ ANTENNA_4/DIODE VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_32_990 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout213_X fanout213/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[0\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1233/X m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/A1 fanout577/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold151 hold151/A VGND VGND VPWR VPWR hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 hold140/A VGND VGND VPWR VPWR hold140/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold162 hold162/A VGND VGND VPWR VPWR hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A VGND VGND VPWR VPWR hold173/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold184 hold184/A VGND VGND VPWR VPWR hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A VGND VGND VPWR VPWR hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout620 fanout621/X VGND VGND VPWR VPWR fanout620/X sky130_fd_sc_hd__buf_2
XFILLER_59_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1 fanout449/X fanout455/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or4_2_A/X fanout444/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1/X sky130_fd_sc_hd__o31a_1
XANTENNA_fanout73_A fanout75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[1\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ hold379/X VGND VGND VPWR VPWR hold378/A sky130_fd_sc_hd__dfxtp_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_4 clkbuf_leaf_19_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4/D
+ VGND VGND VPWR VPWR uo_out[3] sky130_fd_sc_hd__dfxtp_2
XFILLER_73_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__xor2_2_B hold892/A hold767/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
Xdata\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold7/X fanout308/X VGND VGND VPWR VPWR data\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__mux2_1
XFILLER_2_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1003/A fanout56/X fanout28/X m_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.m_matrix\[7\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold980/X hold1027/A fanout545/X VGND VGND VPWR VPWR hold981/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold69/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold93/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[3\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold975/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__xnor2_2_A hold645/A hold376/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout413/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold161/X fanout323/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold855/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A_A m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A0/X hold68/X fanout311/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__a211o_2_A1 hold838/A fanout285/X
+ m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__a22o_2_A1/X fanout372/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_52_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_47_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[5\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[5\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1020/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold292/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_43_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A fanout450/X fanout453/X
+ fanout455/X fanout457/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout194/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A0 hold121/A m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout513/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X m_io.m_config.ll_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold268/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_A2
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A0 hold180/A m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout501/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold752/X hold14/X fanout588/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_B
+ m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_28_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__a211o_2_A1 hold608/A fanout287/X
+ m_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__a22o_2_A1/X fanout396/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A2
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1/Y
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__o311a_4
XPHY_EDGE_ROW_27_Left_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout163_X fanout163/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B/X m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold110/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout330_X fanout330/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/A1
+ fanout104/X ANTENNA_3/DIODE VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_36_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold39/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout402/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[26\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout417/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout450 fanout450/A VGND VGND VPWR VPWR fanout450/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout76_X fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout271/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout461 fanout461/A VGND VGND VPWR VPWR fanout461/X sky130_fd_sc_hd__buf_2
XFILLER_63_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout472 fanout473/X VGND VGND VPWR VPWR fanout472/X sky130_fd_sc_hd__buf_2
XFILLER_48_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout483 fanout484/X VGND VGND VPWR VPWR fanout483/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout494 fanout500/A VGND VGND VPWR VPWR fanout494/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold214/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__and3_2_B_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__a31o_2_A3 fanout446/X fanout479/X
+ hold250/A fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_15_710 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold419/X m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_54_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold41/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_30_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout90 fanout91/A VGND VGND VPWR VPWR fanout90/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A0 hold136/A m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout170/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold909 hold909/A VGND VGND VPWR VPWR hold909/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_B2
+ fanout400/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_A1
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout52/X fanout76/X
+ m_blake2.m_hash256.m_matrix\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21oi_2_A2
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1/X
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2/A1
+ sky130_fd_sc_hd__a21oi_4
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold462/X m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_36_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__inv_2_A hold1212/A VGND VGND VPWR
+ VPWR m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/C
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y_A
+ hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_matrix\[11\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1223/A hold1125/X fanout565/X VGND VGND VPWR VPWR hold1126/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B_A fanout429/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1089/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_80_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout381/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout261/X
+ m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold840/A fanout60/X fanout40/X m_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xnor2_1
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_72_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout351/X m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_20_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold813/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__o31a_2_A3
+ fanout452/X fanout458/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/A
+ sky130_fd_sc_hd__o31a_1
Xm_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold1240/X fanout168/X m_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__nor2_2_B fanout495/X hold166/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__xnor2_2_A hold366/A hold1241/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.g_buffer\[16\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.g_buffer\[11\].m_c_buf m_blake2.m_hash256.g_buffer\[11\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[11\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__a31o_2_A3 fanout446/X fanout478/X
+ hold132/A fanout507/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A_sky130_fd_sc_hd__or2_2_X_B
+ fanout103/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_835 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ hold1244/A fanout357/X fanout269/X m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/B1 sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A0 hold146/A m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A hold467/A m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR ANTENNA_11/DIODE sky130_fd_sc_hd__dfxtp_1
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ fanout612/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2/Y
+ m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout402/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout36_A fanout39/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_B
+ fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1242/A fanout25/X fanout69/X hold662/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_22_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_76_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__xnor2_2_A hold888/A hold685/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_3_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X/C
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout194/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout196/X m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout188/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xfanout280 fanout282/X VGND VGND VPWR VPWR fanout280/X sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_3_Left_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout291 fanout295/A VGND VGND VPWR VPWR fanout291/X sky130_fd_sc_hd__buf_2
XFILLER_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/A1
+ m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/A2 m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/Y sky130_fd_sc_hd__a21oi_1
XFILLER_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold204/X fanout166/X m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_43_871 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold127/X fanout329/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold772/A fanout25/X fanout51/X hold1093/A m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_61_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout153/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout160/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold717 hold717/A VGND VGND VPWR VPWR hold717/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold706 hold706/A VGND VGND VPWR VPWR hold706/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold728 hold728/A VGND VGND VPWR VPWR hold728/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_3_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
Xhold739 hold739/A VGND VGND VPWR VPWR hold739/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout612/X VGND VGND VPWR VPWR m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__and2_1
XFILLER_69_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__a31o_2_B1 hold1008/A
+ m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__and2_2_A/B
+ m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout59/X fanout67/X
+ hold649/A m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A hold502/A hold966/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XFILLER_80_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout240_A fanout240/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A fanout341/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[0\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout126_X fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout505_A fanout509/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__a21oi_2_A1/B1 m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__or2_2
Xm_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/B1
+ sky130_fd_sc_hd__nor2_1
XFILLER_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_1 hold245/A m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout375/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_2
Xm_blake2.m_hash256.m_matrix\[3\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1057/X m_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout588/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y
+ fanout273/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold94/A sky130_fd_sc_hd__dfxtp_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_c_buf\[20\]_sky130_fd_sc_hd__and2_2_X fanout354/X m_blake2.m_hash256.g_c_buf\[20\]_sky130_fd_sc_hd__and2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[20\].m_c_buf/A sky130_fd_sc_hd__and2_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A VGND VGND VPWR VPWR hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A VGND VGND VPWR VPWR hold77/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold88 hold88/A VGND VGND VPWR VPWR hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A VGND VGND VPWR VPWR hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold386/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_3_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold670/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_27_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/B2
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_78_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_8 ANTENNA_8/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[12\].m_y_buf m_blake2.m_hash256.g_buffer\[12\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[12\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_10_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/A1
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/A3
+ m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/X
+ sky130_fd_sc_hd__a32o_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout282/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout195/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold932/X fanout207/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A0 hold928/A m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout523/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/A
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A1 hold381/A m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D
+ sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_50_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_793 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_C
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold1259/A fanout137/X fanout96/X m_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold577/X m_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout597/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1098 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B/Y m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout182/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout156/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold1195/A fanout38/X m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout23/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xhold525 hold525/A VGND VGND VPWR VPWR hold525/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 hold514/A VGND VGND VPWR VPWR hold514/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold536 hold536/A VGND VGND VPWR VPWR hold536/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold503 hold503/A VGND VGND VPWR VPWR hold503/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 hold569/A VGND VGND VPWR VPWR hold569/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and3_2_C_A fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold547 hold547/A VGND VGND VPWR VPWR hold547/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold558 hold558/A VGND VGND VPWR VPWR hold558/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1225 hold1225/A VGND VGND VPWR VPWR hold1225/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout197/X m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout187/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout190_A fanout192/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout229/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1214 hold1214/A VGND VGND VPWR VPWR hold1214/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[13\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[13\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold786/A sky130_fd_sc_hd__dfxtp_1
Xhold1203 hold1203/A VGND VGND VPWR VPWR hold1203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1258 hold1258/A VGND VGND VPWR VPWR hold1258/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__xor2_2_A hold712/A hold807/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_fanout288_A fanout288/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1236 hold1236/A VGND VGND VPWR VPWR hold1236/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1247 hold1247/A VGND VGND VPWR VPWR hold1247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1269 hold794/A VGND VGND VPWR VPWR hold1269/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A1_S fanout323/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__a22o_2_A1 hold644/A fanout289/X
+ fanout285/X hold611/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout243_X fanout243/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold335/A m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout363/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ hold635/X VGND VGND VPWR VPWR hold634/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_22_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__mux2_1_X
+ m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q input14/X fanout1/A VGND VGND VPWR VPWR
+ m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X/B sky130_fd_sc_hd__mux2_1
XANTENNA_fanout410_X fanout410/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A0 hold500/A m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold448/X m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1/X
+ VGND VGND VPWR VPWR fanout232/A sky130_fd_sc_hd__and2b_4
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold783/X m_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout549/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1 hold235/A fanout102/X
+ m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1/B1 m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A1 sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold533/X m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1227/A fanout81/X fanout73/X m_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_5_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_B1
+ fanout346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout349/X m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a21o_1
XFILLER_45_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__or2_2_B fanout488/X hold151/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__a22o_2_A1 hold342/A fanout190/X
+ fanout198/X hold964/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/A2
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_73_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_13_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B fanout452/X fanout454/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_2
Xm_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ hash\[6\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold715/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_A2 m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold955/X hold1031/X fanout592/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/A1
+ m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/A2 m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/X sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_52_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout278/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1062/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout583/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/A fanout220/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XFILLER_35_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold740/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout413/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout520/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__mux2_1_A1_S fanout208/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1/B2
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_52_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold30/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold337/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[31\]_sky130_fd_sc_hd__or2_2_A hold538/A fanout392/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[31\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[13\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1024/A sky130_fd_sc_hd__dfxtp_1
Xhold311 hold311/A VGND VGND VPWR VPWR hold311/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold300 hold300/A VGND VGND VPWR VPWR hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold322 hold322/A VGND VGND VPWR VPWR hold322/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout203_A fanout204/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold344 hold344/A VGND VGND VPWR VPWR hold344/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 hold333/A VGND VGND VPWR VPWR hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold366 hold366/A VGND VGND VPWR VPWR hold366/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 hold377/A VGND VGND VPWR VPWR hold377/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[1\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[1\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold947/A sky130_fd_sc_hd__dfxtp_1
Xhold355 hold355/A VGND VGND VPWR VPWR hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold399 hold399/A VGND VGND VPWR VPWR hold399/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold391/X fanout207/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold432/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold678/X m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold388 hold388/A VGND VGND VPWR VPWR hold388/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input8_A ui_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 hold1000/A VGND VGND VPWR VPWR hold1000/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout193_X fanout193/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1022 hold1022/A VGND VGND VPWR VPWR hold1022/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1033 hold1033/A VGND VGND VPWR VPWR hold1033/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_24_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1011 hold1011/A VGND VGND VPWR VPWR hold1011/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1127/A sky130_fd_sc_hd__dfxtp_1
Xhold1055 hold1055/A VGND VGND VPWR VPWR hold1055/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1066 hold1066/A VGND VGND VPWR VPWR hold1066/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1044 hold1044/A VGND VGND VPWR VPWR hold1044/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 hold1088/A VGND VGND VPWR VPWR hold1088/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1099 hold1099/A VGND VGND VPWR VPWR hold1099/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_c_buf\[12\]_sky130_fd_sc_hd__a211o_2_X hold793/A fanout174/X
+ m_blake2.m_hash256.g_c_buf\[12\]_sky130_fd_sc_hd__a211o_2_X/B1 m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__a32o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[12\].m_c_buf/A sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__and2_2_B_A fanout429/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1077 hold1077/A VGND VGND VPWR VPWR hold1077/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold532/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A fanout219/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout285/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold926/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold92/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__and3_2_A hold213/A fanout463/X fanout368/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold567/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold442/X m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold804/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold368/X fanout335/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__a22o_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_43_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold539/X hold995/A fanout600/X VGND VGND VPWR VPWR hold540/A sky130_fd_sc_hd__mux2_1
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold545/X m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout160/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1129/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__or2_2_A hold1235/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout268/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.g_buffer\[18\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_58_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B fanout490/X hold120/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_79_1430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__o21a_2_A1 m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/A
+ fanout379/X fanout407/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_17_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_955 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_15_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_2
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_45_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[12\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1210/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_41_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold864/A m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout502/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1238/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold675/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold301/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[12\]\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1244/X fanout228/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1236/X m_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout566/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_idx_next\[0\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B fanout481/X VGND
+ VGND VPWR VPWR fanout303/A sky130_fd_sc_hd__and3_2
Xfanout109 fanout111/A VGND VGND VPWR VPWR fanout109/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__inv_2_A fanout495/X VGND VGND VPWR
+ VPWR fanout443/A sky130_fd_sc_hd__inv_2
Xm_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/X fanout609/X input3/X VGND VGND VPWR VPWR m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[14\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold538/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout153/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold296/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[2\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ hold728/X VGND VGND VPWR VPWR hold727/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout153_A fanout154/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_2
XFILLER_1_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__a221o_2_A1 hold1174/A fanout276/X
+ fanout176/A m_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__or2_2_A/X fanout272/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout320_A fanout323/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__o2bb2a_2_A1_N hold390/A fanout304/X fanout374/X
+ hold907/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X
+ sky130_fd_sc_hd__o2bb2a_1
Xm_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold298/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__inv_2_Y
+ fanout469/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ sky130_fd_sc_hd__inv_6
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_30_clk clkload4/A VGND VGND VPWR VPWR clkbuf_leaf_30_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout418_A fanout420/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A1_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__and3_2_C fanout447/X fanout480/X
+ hold145/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2 m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ fanout261/X fanout306/X m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__or2_2_A/A VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/X sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__or2_2_A hold281/A fanout364/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhold152 hold152/A VGND VGND VPWR VPWR hold152/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 hold130/A VGND VGND VPWR VPWR hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 hold141/A VGND VGND VPWR VPWR hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/A VGND VGND VPWR VPWR hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/A VGND VGND VPWR VPWR hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[4\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold958/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[8\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold819/A sky130_fd_sc_hd__dfxtp_1
Xhold163 hold163/A VGND VGND VPWR VPWR hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout610 fanout615/X VGND VGND VPWR VPWR fanout610/X sky130_fd_sc_hd__clkbuf_2
Xfanout621 input2/X VGND VGND VPWR VPWR fanout621/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold196 hold196/A VGND VGND VPWR VPWR hold196/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__nor2_2_B fanout483/X hold106/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1230/X fanout223/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_S fanout218/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_5 clkbuf_leaf_19_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5/D
+ VGND VGND VPWR VPWR uo_out[2] sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[6\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[6\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1033/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_928 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout444/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/X m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_21_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkload15/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold37/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__a211oi_2_A1 hold411/A fanout288/X
+ m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__a22o_2_A1/X fanout378/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__a211oi_2_A1/Y
+ sky130_fd_sc_hd__a211oi_1
Xm_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold498/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout259/X m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR fanout176/A sky130_fd_sc_hd__nor2_4
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[8\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold577/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__a21o_2_X
+ fanout284/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_A1/Y fanout466/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X/C
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_34_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X hold1162/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[29\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__xor2_2_A hold262/A hold591/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold87/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A2 m_io.cmd\[5\]_sky130_fd_sc_hd__and2b_2_B/X
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_72_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1093/A fanout99/X fanout148/X hold503/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_43_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold960/A sky130_fd_sc_hd__dfxtp_1
Xdata_idx\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X hold5/X VGND VGND VPWR
+ VPWR data_idx\[0\]_sky130_fd_sc_hd__and4_2_B/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold121/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__nand2_2_B fanout431/X hold175/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ hold765/X VGND VGND VPWR VPWR hold764/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_12_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_12_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold180/X fanout310/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout188/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout196/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__mux2_1_A1_S fanout341/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout200/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A hold357/A fanout288/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_68_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A1_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout270_A fanout271/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A0_S fanout520/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ hold670/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__o21a_2_A1 hold776/A fanout366/X
+ fanout169/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[8\]_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout156_X fanout156/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ sky130_fd_sc_hd__a21oi_2
XANTENNA_data\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A0 hold66/A m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold849/X hold1096/A fanout555/X VGND VGND VPWR VPWR hold850/A sky130_fd_sc_hd__mux2_1
XFILLER_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout323_X fanout323/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold393/X m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__xnor2_2_A hold832/A hold682/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout300/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout440 fanout441/X VGND VGND VPWR VPWR fanout440/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout176/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout451 fanout453/X VGND VGND VPWR VPWR fanout451/X sky130_fd_sc_hd__buf_2
XFILLER_63_1072 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout462 hold1180/A VGND VGND VPWR VPWR fanout462/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold107/A sky130_fd_sc_hd__dfxtp_1
Xfanout473 fanout473/A VGND VGND VPWR VPWR fanout473/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold191/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xfanout484 fanout486/X VGND VGND VPWR VPWR fanout484/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_matrix\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold988/X hold967/X fanout584/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout495 fanout497/X VGND VGND VPWR VPWR fanout495/X sky130_fd_sc_hd__clkbuf_4
Xm_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ hold6/A m_io.data_v_early_sky130_fd_sc_hd__and3_2_C/X hold2/X VGND VGND VPWR VPWR
+ m_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y/B
+ sky130_fd_sc_hd__a21oi_1
XFILLER_59_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold202/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_30_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1119/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold893/X hold435/X fanout558/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout91 fanout91/A VGND VGND VPWR VPWR fanout91/X sky130_fd_sc_hd__buf_2
XFILLER_31_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout80 fanout83/A VGND VGND VPWR VPWR fanout80/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold136/X fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xor2_4
XFILLER_35_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold656/A fanout55/X fanout42/X m_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__xnor2_2_A hold272/A m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2/X
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.m_matrix\[7\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold606/X hold1179/A fanout588/X VGND VGND VPWR VPWR hold607/A sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_1_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_1_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X m_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold218/A sky130_fd_sc_hd__dfxtp_1
XFILLER_64_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A0 hold32/A m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_S fanout214/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/A
+ m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2 hold514/A m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/D
+ sky130_fd_sc_hd__and4_2
Xm_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__xnor2_2_A hold420/A hold226/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout157/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_S fanout415/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_A fanout119/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__xnor2_2_B hold760/A hold838/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold789/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout485_A fanout486/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold89/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold780/A fanout109/X fanout121/X hold1201/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_buffer\[15\].m_c_buf m_blake2.m_hash256.g_buffer\[15\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[15\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/A1
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/X
+ sky130_fd_sc_hd__o21ba_1
XFILLER_18_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A/A
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_56_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout273_X fanout273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_858 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_880 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold146/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__o21bai_2_A1/Y m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/X
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__nand3_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_X fanout538/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/D
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ sky130_fd_sc_hd__a21o_1
XFILLER_12_703 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout181/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_C
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_A fanout408/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A2
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_matrix\[5\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold768/X hold700/X fanout553/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xclkload0 clkload0/A VGND VGND VPWR VPWR clkload0/Y sky130_fd_sc_hd__bufinv_16
XTAP_TAPCELL_ROW_22_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_c_buf\[8\]_sky130_fd_sc_hd__a211o_2_X hold730/A fanout174/X
+ m_blake2.m_hash256.g_c_buf\[8\]_sky130_fd_sc_hd__a211o_2_X/B1 m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__a32o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[8\].m_c_buf/A sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_76_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_72_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.g_buffer\[22\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[1\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout209/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_43_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout270 fanout271/X VGND VGND VPWR VPWR fanout270/X sky130_fd_sc_hd__clkbuf_4
XFILLER_43_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout281 fanout282/X VGND VGND VPWR VPWR fanout281/X sky130_fd_sc_hd__clkbuf_2
Xfanout292 fanout294/X VGND VGND VPWR VPWR fanout292/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[3\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ hold882/X VGND VGND VPWR VPWR hold881/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_B2
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A0 hold154/A m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout181/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_S fanout203/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1238/A fanout50/X fanout38/X hold582/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout128/X
+ fanout112/X hold918/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ hold21/X m_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/A2
+ fanout611/X VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xhash\[3\]_sky130_fd_sc_hd__mux2_1_A0 hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout485/X VGND VGND VPWR VPWR hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_4
XTAP_TAPCELL_ROW_61_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[0\].m_y_buf m_blake2.m_hash256.g_buffer\[0\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[0\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__xor2_2_B hold323/A hold761/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A fanout152/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ hold1075/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xhold718 hold718/A VGND VGND VPWR VPWR hold718/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_S fanout418/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold707 hold707/A VGND VGND VPWR VPWR hold707/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold729 hold729/A VGND VGND VPWR VPWR hold729/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__xnor2_2_A hold855/A hold800/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold658/X hold1117/A fanout580/X VGND VGND VPWR VPWR hold659/A sky130_fd_sc_hd__mux2_1
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout417/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__or2_2_A hold390/X fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout89/X m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/B1
+ sky130_fd_sc_hd__a211o_1
XFILLER_78_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1056/A fanout70/X fanout74/X hold967/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__and3_2_B_B
+ m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.f_finished_q_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X/A1
+ m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X/A2 m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR ANTENNA_4/DIODE sky130_fd_sc_hd__o21a_1
XFILLER_37_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a31o_2_X
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0_S fanout299/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X
+ fanout119/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__xnor2_2_A hold418/A hold618/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_B1
+ fanout354/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout233_A fanout234/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold340/X m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/B m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A/X
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a221o_2_C1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout400_A fanout400/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A/A
+ m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold315/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ fanout239/X m_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A/C
+ sky130_fd_sc_hd__inv_2
XFILLER_9_1370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_57_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold89 hold89/A VGND VGND VPWR VPWR hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A VGND VGND VPWR VPWR hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A VGND VGND VPWR VPWR hold78/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__or2_2_A_B fanout243/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout53/X
+ fanout37/X hold1085/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold364/X
+ fanout161/X m_io.m_config.ll_q\[9\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_45_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[22\]_sky130_fd_sc_hd__mux2_1_A1_S fanout223/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_S fanout231/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_9 fanout43/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhash_v_sky130_fd_sc_hd__a211o_2_X fanout463/X hash_v_sky130_fd_sc_hd__a211o_2_X/A2
+ hold21/X fanout478/X VGND VGND VPWR VPWR hash_v_sky130_fd_sc_hd__a211o_2_X/X sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[16\].m_y_buf m_blake2.m_hash256.g_buffer\[16\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[16\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold145/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold289/X fanout167/X m_io.m_config.ll_q\[12\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_66_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y
+ fanout83/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_B1 fanout100/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold928/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__xnor2_2_B hold1214/A hold754/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o21a_2_A2
+ fanout452/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_16_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_0_clk_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__mux2_1_A0 hold270/A m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout371/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/A2
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X fanout402/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1
+ fanout400/X m_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout267/X m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1/X
+ sky130_fd_sc_hd__o221a_1
Xhold526 hold526/A VGND VGND VPWR VPWR hold526/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_B1_sky130_fd_sc_hd__or3_2_X
+ fanout407/X fanout458/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2/B1
+ sky130_fd_sc_hd__or3_1
XANTENNA_m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold515 hold515/A VGND VGND VPWR VPWR hold515/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold504 hold504/A VGND VGND VPWR VPWR hold504/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and3_2_C_B fanout478/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
Xhold548 hold548/A VGND VGND VPWR VPWR hold548/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold537 hold537/A VGND VGND VPWR VPWR hold537/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 hold559/A VGND VGND VPWR VPWR hold559/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nor2_1
Xhold1215 hold1215/A VGND VGND VPWR VPWR hold1215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1204 hold1204/A VGND VGND VPWR VPWR hold1204/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1226 hold1226/A VGND VGND VPWR VPWR hold1226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1237 hold1237/A VGND VGND VPWR VPWR hold1237/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1248 hold1248/A VGND VGND VPWR VPWR hold1248/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ fanout169/X m_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout251/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout183_A fanout184/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1259 hold1259/A VGND VGND VPWR VPWR hold1259/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_0_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout350_A fanout361/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__xnor2_2_A hold905/A hold465/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold279/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold752/A fanout62/X fanout42/X m_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold995/A fanout131/X fanout147/X hold630/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_24_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X hold483/A fanout18/X m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[26\].m_y_buf/A sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout615_A input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold335/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout236_X fanout236/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold1029/A fanout116/X fanout99/X hold722/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold17/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold614/X fanout164/X m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__or2_2_A/X fanout617/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout160/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold323/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout403_X fanout403/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout559/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__or2_2_B_A fanout494/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout300/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold500/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1014/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout96_A fanout99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_735 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__nand2_2_B fanout439/X hold170/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y/A2
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold821/A fanout111/X fanout114/X hold1195/A m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A/X fanout611/X VGND VGND VPWR VPWR
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1
+ fanout400/X m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout266/X fanout366/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA_clkbuf_leaf_2_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold603/X m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout212/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1234/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[12\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold319/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
XFILLER_32_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold251/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold492/A m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout372/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B fanout484/X hold288/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A
+ fanout170/X fanout172/X m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A2
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A_B m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__and2_2_A/X sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout186/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_X
+ fanout249/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_1 hold221/A m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout397/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold85/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/C
+ sky130_fd_sc_hd__nand2_1
XFILLER_80_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout422/A m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1/B1
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold588/X m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout413/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_35_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_A1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_B2
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold191/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__or2_2_B_A fanout497/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__nor2_2_B_A fanout478/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold57/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout178/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold254/X m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold301 hold301/A VGND VGND VPWR VPWR hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout414/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold618/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold312 hold312/A VGND VGND VPWR VPWR hold312/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X
+ hold1219/A fanout393/X fanout239/X m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/A1 sky130_fd_sc_hd__o211a_1
Xhold334 hold334/A VGND VGND VPWR VPWR hold334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 hold323/A VGND VGND VPWR VPWR hold323/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout125/X
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a21o_1
Xhold378 hold378/A VGND VGND VPWR VPWR hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 hold356/A VGND VGND VPWR VPWR hold356/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold345 hold345/A VGND VGND VPWR VPWR hold345/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 hold367/A VGND VGND VPWR VPWR hold367/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold389 hold389/A VGND VGND VPWR VPWR hold389/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C_A
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_A fanout399/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X
+ hold700/A fanout112/X fanout116/X m_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A3
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_5_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1001 hold1001/A VGND VGND VPWR VPWR hold1001/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1023 hold1023/A VGND VGND VPWR VPWR hold1023/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[1\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold553/X hold1192/A fanout556/X VGND VGND VPWR VPWR hold554/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1078/A fanout84/X fanout136/X hold920/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xhold1012 hold1012/A VGND VGND VPWR VPWR hold1012/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 hold1067/A VGND VGND VPWR VPWR hold1067/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 hold1056/A VGND VGND VPWR VPWR hold1056/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout186_X fanout186/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1034 hold1034/A VGND VGND VPWR VPWR hold1034/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_2
XFILLER_39_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1045 hold1045/A VGND VGND VPWR VPWR hold1045/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold320/A m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout375/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout258/X m_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout383/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
Xhold1089 hold1089/A VGND VGND VPWR VPWR hold1089/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1078 hold1078/A VGND VGND VPWR VPWR hold1078/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold596/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold790/A fanout131/X fanout99/X hold992/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__o21a_2_A1 hold916/A fanout362/X
+ fanout171/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_14_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout520_X fanout520/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3_2_B/A
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A0 hold129/A m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A_A m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout184/X m_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_B_A_N
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_A
+ fanout269/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1192/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
Xm_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__or4_2_B hold6/A hold3/A hold4/A
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__or4_2_B/D VGND VGND VPWR VPWR
+ block_last_sky130_fd_sc_hd__a32o_2_B2/B1 sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold374/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout184/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_2
XFILLER_27_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold890 hold890/A VGND VGND VPWR VPWR hold890/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A/Y m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout260/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1/X
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ sky130_fd_sc_hd__a31o_1
XFILLER_79_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A_B m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ fanout487/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_72_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[3\]_sky130_fd_sc_hd__mux2_1_A0 hold1185/X m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout236/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold699/X VGND VGND VPWR VPWR hold698/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1069/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_hash\[3\]_sky130_fd_sc_hd__mux2_1_A0_S fanout485/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_4
Xm_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold972/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold911/X hold820/X fanout597/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold864/X fanout309/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_S fanout419/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold847/A fanout130/X fanout134/X hold924/A m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__a21oi_2_B1_B1 m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_B2_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1/B2 sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold40/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold550/X m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[5\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1195/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold463/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__nor2_2_B fanout478/X hold185/A VGND
+ VGND VPWR VPWR fanout427/A sky130_fd_sc_hd__nor2_1
XFILLER_67_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.g_buffer\[24\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_io.m_block_data.data_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ hold6/A m_io.data_v_early_sky130_fd_sc_hd__and3_2_C/X m_io.m_block_data.data_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A0 hold113/A m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[1\]_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__or3b_2_X
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/A m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[1\]_sky130_fd_sc_hd__and2b_2_X/B
+ sky130_fd_sc_hd__or3b_1
XFILLER_36_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X m_io.m_config.ll_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold364/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/D
+ m_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xm_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__or2_2_A hold334/A fanout248/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_51_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__a22o_2_A1 hold843/A fanout280/X
+ fanout287/X hold653/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A0 hold184/A m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold183/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold865/A fanout26/X fanout54/X hold1187/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout146_A fanout147/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/B m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/D
+ sky130_fd_sc_hd__and4_1
XFILLER_52_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1208/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold48/A m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout529/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout313_A fanout314/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout485/X VGND VGND VPWR VPWR m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xhold142 hold142/A VGND VGND VPWR VPWR hold142/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A VGND VGND VPWR VPWR hold131/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold153 hold153/A VGND VGND VPWR VPWR hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold120/A VGND VGND VPWR VPWR hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A VGND VGND VPWR VPWR hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A VGND VGND VPWR VPWR hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A VGND VGND VPWR VPWR hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 fanout612/X VGND VGND VPWR VPWR fanout611/X sky130_fd_sc_hd__buf_2
Xfanout600 fanout602/X VGND VGND VPWR VPWR fanout600/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/A2
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__and2b_2
Xm_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__or2_2_A hold1166/A fanout362/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_8_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold197 hold197/A VGND VGND VPWR VPWR hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[10\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1187/X m_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout593/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[4\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1108/X hold1079/X fanout555/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_6 clkbuf_leaf_19_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6/D
+ VGND VGND VPWR VPWR uo_out[1] sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1
+ fanout375/X m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1/X fanout188/X fanout178/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2/B1
+ sky130_fd_sc_hd__a221o_1
XFILLER_54_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_1047 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_992 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A_B
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout231/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__a22o_2_A1 hold437/X fanout319/X
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__a22o_2_A1/B1 fanout512/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold326/A m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__and2_2_B/X fanout376/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[4\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold943/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_9_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_B2
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout48/X fanout36/X
+ hold1020/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_34_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout514/X m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_34_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y/A m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A0 hold229/A m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout501/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_47_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_47_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout232/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[12\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold952/A hold424/X fanout586/X VGND VGND VPWR VPWR hold425/A sky130_fd_sc_hd__mux2_1
XFILLER_9_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__inv_2_A m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.m_matrix\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold747/X hold680/X fanout576/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1188/X m_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout540/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold694/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1111/X hold1093/X fanout573/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__and3_2_A hold201/A fanout465/X fanout395/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1 hold1128/A fanout347/X
+ fanout260/X m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/B2 fanout268/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1190/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_42_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2
+ fanout240/X m_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__or2_2_A/A m_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XANTENNA_fanout430_A fanout431/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold926/A fanout82/X fanout70/X hold601/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold66/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout153/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold1236/A fanout53/X fanout81/X m_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__xnor2_2_A hold623/A hold932/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__and2_2_B fanout439/X hold90/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[5\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold530/A fanout90/X fanout130/X hold577/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_48_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout430 fanout431/X VGND VGND VPWR VPWR fanout430/X sky130_fd_sc_hd__clkbuf_4
Xfanout441 fanout442/X VGND VGND VPWR VPWR fanout441/X sky130_fd_sc_hd__clkbuf_4
Xfanout463 fanout465/A VGND VGND VPWR VPWR fanout463/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__xnor2_2_A hold446/A hold737/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xfanout452 fanout453/X VGND VGND VPWR VPWR fanout452/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout474 fanout475/X VGND VGND VPWR VPWR fanout474/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.g_buffer\[3\].m_c_buf m_blake2.m_hash256.g_buffer\[3\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[3\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout485 fanout486/X VGND VGND VPWR VPWR fanout485/X sky130_fd_sc_hd__clkbuf_4
Xfanout496 fanout497/X VGND VGND VPWR VPWR fanout496/X sky130_fd_sc_hd__buf_2
XANTENNA_m_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__or2_2_A_B fanout248/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/A1
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/A2
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/A3
+ fanout104/X m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__a32o_4
XFILLER_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__o21ai_2_A1 hold560/A fanout375/X
+ fanout193/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_30_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout70 fanout71/A VGND VGND VPWR VPWR fanout70/X sky130_fd_sc_hd__clkbuf_4
Xfanout92 fanout95/A VGND VGND VPWR VPWR fanout92/X sky130_fd_sc_hd__buf_4
Xfanout81 fanout83/A VGND VGND VPWR VPWR fanout81/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__xnor2_2_A hold804/A hold806/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XFILLER_10_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_36_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_A2_sky130_fd_sc_hd__or4_2_X
+ fanout455/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/C m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/A2
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold632/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1_S fanout218/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold32/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.res_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XFILLER_33_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1384 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__and2_2_A/B fanout423/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XANTENNA_m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B_A fanout499/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[15\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold720/X hold549/X fanout560/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout109_A fanout111/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A hold256/A m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout351/X m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__a22o_2_A1/X fanout180/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A fanout480/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X m_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold605/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
XFILLER_25_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A0 hold27/A m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout266_X fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_buffer\[19\].m_c_buf m_blake2.m_hash256.g_buffer\[19\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[19\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2 m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ fanout260/X fanout305/X m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/C1
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/X sky130_fd_sc_hd__a221o_1
XFILLER_52_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__nand2_2_B/Y
+ fanout266/X fanout389/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_34_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__xnor2_2_A hold298/A hold387/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_715 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload1 clkload1/A VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__inv_6
XFILLER_32_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_76_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold672/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold155/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold796/A sky130_fd_sc_hd__dfxtp_1
Xfanout260 fanout265/X VGND VGND VPWR VPWR fanout260/X sky130_fd_sc_hd__clkbuf_4
Xfanout271 fanout273/A VGND VGND VPWR VPWR fanout271/X sky130_fd_sc_hd__clkbuf_4
Xfanout282 fanout283/X VGND VGND VPWR VPWR fanout282/X sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold730/X fanout221/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout293 fanout294/X VGND VGND VPWR VPWR fanout293/X sky130_fd_sc_hd__buf_2
XFILLER_74_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N/Y
+ sky130_fd_sc_hd__o21bai_2
Xm_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold154/X fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__nand2_2_B fanout438/X hold205/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X hash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_851 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__o21a_2_A1 hold743/A fanout366/X
+ fanout250/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold336/X m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ fanout160/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N/X
+ sky130_fd_sc_hd__o21ba_1
Xm_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout255/X m_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ fanout369/X fanout177/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_61_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout117/X
+ fanout145/X m_blake2.m_hash256.m_matrix\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
Xhold708 hold708/A VGND VGND VPWR VPWR hold708/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout181/X m_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_2
Xhold719 hold719/A VGND VGND VPWR VPWR hold719/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold499/X m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X fanout413/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[4\].m_y_buf m_blake2.m_hash256.g_buffer\[4\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[4\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A0 hold101/A m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout280/X m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ hold1052/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 fanout240/X hold1064/A
+ m_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XFILLER_38_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B_A fanout489/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold914/X m_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout593/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A0 hold158/A m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ fanout237/X m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
XFILLER_37_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_A1
+ fanout288/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout345/X m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__nor2_1
XFILLER_34_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2_B1 fanout307/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_A fanout228/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold508/X hold351/X fanout560/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__or2_2_B fanout493/X hold215/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_20_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_906 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout195/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_60_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A VGND VGND VPWR VPWR hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_25_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold68 hold68/A VGND VGND VPWR VPWR hold68/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_buffer\[30\].m_c_buf m_blake2.m_hash256.g_buffer\[30\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[30\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_854 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XFILLER_40_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C/X
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/B
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__a31o_2_A3 fanout448/X fanout480/X
+ hold181/A fanout534/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.g_c_buf\[30\]_sky130_fd_sc_hd__a22o_2_X fanout355/X m_blake2.m_hash256.g_c_buf\[30\]_sky130_fd_sc_hd__a22o_2_X/A2
+ m_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__or2_2_A/X fanout253/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[30\].m_c_buf/A sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__nand2_1
XFILLER_10_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_A
+ fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/X
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/A
+ sky130_fd_sc_hd__a21o_2
XFILLER_3_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold1115/A fanout86/X fanout98/X hold1033/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_63_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkload4_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold638/X hold930/A fanout588/X VGND VGND VPWR VPWR hold639/A sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ fanout451/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
XFILLER_37_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2/B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_71_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold313/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_50_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand3_2_B
+ m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/C
+ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_13_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y/A
+ sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1
+ fanout288/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout295/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold505 hold505/A VGND VGND VPWR VPWR hold505/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 hold516/A VGND VGND VPWR VPWR hold516/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 hold527/A VGND VGND VPWR VPWR hold527/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1 hold525/A fanout256/X
+ fanout196/X hold593/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xhold538 hold538/A VGND VGND VPWR VPWR hold538/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 hold549/A VGND VGND VPWR VPWR hold549/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1194/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_X
+ m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold1216 hold1216/A VGND VGND VPWR VPWR hold1216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1205 hold1205/A VGND VGND VPWR VPWR hold1205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1238 hold1238/A VGND VGND VPWR VPWR hold1238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1249 hold1249/A VGND VGND VPWR VPWR hold1249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1227 hold1227/A VGND VGND VPWR VPWR hold1227/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_69_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[12\]\[2\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold997/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout176_A fanout176/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold685/X m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout299/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__or2_2_A hold218/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold959/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout229_X fanout229/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A
+ hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold711/X m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold851/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold937/X m_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout557/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ fanout452/X fanout152/X m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout482/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ hold1083/A fanout349/X fanout268/X m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__a22o_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X/B1 sky130_fd_sc_hd__a211o_1
XFILLER_49_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold551/A fanout48/X fanout68/X m_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1156/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[15\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1201/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold731/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold504/X m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout44_X fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold458/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_24_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold492/X fanout410/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1007/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A ANTENNA_8/DIODE m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold438/X m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout123/X
+ fanout150/X m_blake2.m_hash256.m_matrix\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold406/X m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_56_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__o21a_2_A1 hold1030/A fanout388/X
+ fanout408/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold506/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_block_data.data_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_io.m_block_data.data_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold4/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_56_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout160/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[31\].m_y_buf m_blake2.m_hash256.g_buffer\[31\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[31\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_43_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[11\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold732/X m_blake2.m_hash256.m_matrix\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout586/X
+ VGND VGND VPWR VPWR hold733/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout290/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y/B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_78_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1/Y sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[8\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold407/X m_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout540/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_B
+ m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold283/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold413/A m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout389/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A1_S fanout411/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout409/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A1
+ fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N_A_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold461/X
+ fanout165/X m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xhold302 hold302/A VGND VGND VPWR VPWR hold302/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 hold313/A VGND VGND VPWR VPWR hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 hold324/A VGND VGND VPWR VPWR hold324/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 hold335/A VGND VGND VPWR VPWR hold335/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xhold368 hold368/A VGND VGND VPWR VPWR hold368/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 hold346/A VGND VGND VPWR VPWR hold346/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 hold357/A VGND VGND VPWR VPWR hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold379 hold379/A VGND VGND VPWR VPWR hold379/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold347/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1270/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout293_A fanout294/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1024 hold1024/A VGND VGND VPWR VPWR hold1024/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1/B1
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold562/X m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 hold1013/A VGND VGND VPWR VPWR hold1013/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1002 hold1002/A VGND VGND VPWR VPWR hold1002/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1057 hold1057/A VGND VGND VPWR VPWR hold1057/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold998/A fanout110/X fanout130/X hold646/A m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xhold1046 hold1046/A VGND VGND VPWR VPWR hold1046/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 hold1035/A VGND VGND VPWR VPWR hold1035/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold320/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold1068 hold1068/A VGND VGND VPWR VPWR hold1068/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout179_X fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1079 hold1079/A VGND VGND VPWR VPWR hold1079/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout291/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold329/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold1143/X fanout162/X m_io.m_config.ll_q\[10\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X
+ VGND VGND VPWR VPWR hold1144/A sky130_fd_sc_hd__o211a_1
XANTENNA_fanout346_X fanout346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold783/A fanout48/X m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__a22o_2_A1 hold97/X fanout317/X
+ m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__a22o_2_A1/B1 fanout508/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold129/X fanout340/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold933/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold444/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A/A
+ fanout320/X m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[8\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1191/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.v_q\[8\]\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold951/X fanout224/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1_Y m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold891 hold891/A VGND VGND VPWR VPWR hold891/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout288/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold880 hold880/A VGND VGND VPWR VPWR hold880/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__and2_2_B_A fanout430/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2
+ fanout260/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout118/X
+ fanout98/X hold1238/A m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold628/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_blake2.m_hash256.round_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout456/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2/X
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XFILLER_13_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1006/X fanout576/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_S fanout303/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1090/X hold1039/X fanout578/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[1\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1242/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X/B
+ sky130_fd_sc_hd__nand3_1
XFILLER_4_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold1204/A fanout57/X fanout25/X hold1041/A m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1202/A fanout24/X fanout32/X m_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold213/X fanout161/X m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__or2_2_A/X fanout614/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_80_1057 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold119/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold116/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_idx\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X hold3/X VGND VGND VPWR
+ VPWR data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/C sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold113/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold771/X fanout554/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__nand2_2_B_A fanout431/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_732 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X
+ hold909/A fanout101/X m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B/A
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ fanout359/X m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X fanout257/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_36_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold184/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A hold437/A VGND VGND VPWR
+ VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_24_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold200/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XFILLER_50_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold627/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold712/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold48/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout306_A fanout307/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ hold891/X VGND VGND VPWR VPWR hold890/A sky130_fd_sc_hd__dfxtp_1
Xhold110 hold110/A VGND VGND VPWR VPWR hold110/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 hold121/A VGND VGND VPWR VPWR hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 hold132/A VGND VGND VPWR VPWR hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout182/X m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_4
Xhold143 hold143/A VGND VGND VPWR VPWR hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold165 hold165/A VGND VGND VPWR VPWR hold165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 hold176/A VGND VGND VPWR VPWR hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 hold154/A VGND VGND VPWR VPWR hold154/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout612 fanout615/X VGND VGND VPWR VPWR fanout612/X sky130_fd_sc_hd__buf_2
XFILLER_63_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout601 fanout602/X VGND VGND VPWR VPWR fanout601/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold187 hold187/A VGND VGND VPWR VPWR hold187/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold198 hold198/A VGND VGND VPWR VPWR hold198/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_S fanout208/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_X fanout296/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A1
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1228/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1_S fanout377/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout100/X hold508/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o32a_2
Xm_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold116/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_buffer\[30\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A0 hold203/A m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout463_X fanout463/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.ll_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold371/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__o21a_2_A1 hold721/A fanout365/X
+ fanout250/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_2_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_7 clkbuf_leaf_20_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7/D
+ VGND VGND VPWR VPWR uo_out[0] sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_S fanout215/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A0 hold443/A m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_1059 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold939/A fanout89/X fanout141/X hold1242/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1155/A fanout29/X fanout65/X hold1063/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__xnor2_2_A hold335/A hold837/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_30_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__nor2_4
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_70_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__a221o_2_B2 hold965/A fanout352/X fanout307/X
+ hold289/A fanout269/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__a221o_2_B2/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_S fanout414/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_9_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X
+ hold786/A fanout30/X fanout82/X hold1103/A m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_34_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR ANTENNA_5/DIODE sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_34_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold229/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_47_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout63/X
+ fanout83/X hold319/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X_B1 m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold403/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout100/X hold894/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o32a_2
Xm_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold213/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A hold478/A m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B fanout489/X ANTENNA_5/DIODE
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout192/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout101/X m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/A1 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/A
+ sky130_fd_sc_hd__o32a_4
XFILLER_68_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__a211o_2_A1 hold466/A fanout280/X
+ m_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__a22o_2_A1/X fanout389/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A0 hold183/A m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/D
+ m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1085/A fanout112/X fanout141/X m_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_64_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout256_A fanout258/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout102/X hold453/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o32a_2
XFILLER_24_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_908 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout211_X fanout211/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_S fanout420/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__and2_2_B_A fanout442/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout431 fanout443/X VGND VGND VPWR VPWR fanout431/X sky130_fd_sc_hd__buf_2
Xfanout420 fanout420/A VGND VGND VPWR VPWR fanout420/X sky130_fd_sc_hd__buf_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout275/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout464 fanout465/X VGND VGND VPWR VPWR fanout464/X sky130_fd_sc_hd__buf_2
Xfanout453 fanout453/A VGND VGND VPWR VPWR fanout453/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout475 fanout476/X VGND VGND VPWR VPWR fanout475/X sky130_fd_sc_hd__buf_4
XANTENNA_fanout71_A fanout71/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout442 fanout443/X VGND VGND VPWR VPWR fanout442/X sky130_fd_sc_hd__clkbuf_4
Xfanout486 fanout500/A VGND VGND VPWR VPWR fanout486/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_59_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout497 fanout500/X VGND VGND VPWR VPWR fanout497/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[7\].m_c_buf m_blake2.m_hash256.g_buffer\[7\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[7\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y fanout273/X m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_27_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout55/X
+ fanout35/X m_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout71 fanout71/A VGND VGND VPWR VPWR fanout71/X sky130_fd_sc_hd__clkbuf_2
Xfanout82 fanout83/A VGND VGND VPWR VPWR fanout82/X sky130_fd_sc_hd__clkbuf_4
Xfanout60 fanout63/X VGND VGND VPWR VPWR fanout60/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout93 fanout95/A VGND VGND VPWR VPWR fanout93/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__mux2_1_A0 hold717/X m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/B1 m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B/C
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.g_buffer\[27\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Left_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout446/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold668/X hold974/A fanout601/X VGND VGND VPWR VPWR hold669/A sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1050/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A0 hold249/A m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout502/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__xnor2_2_A hold545/A hold285/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__or2_2_A hold223/A fanout369/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__a21oi_2_B1 m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ hash\[2\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_32_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2
+ fanout354/X m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_20_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__mux2_1_A1_S fanout228/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_S fanout223/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_21_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1 hold859/A fanout388/X
+ fanout249/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_14_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__xnor2_2_A hold972/A hold578/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B_B m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout231/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_41_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout237/X m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
Xclkload30 clkload30/A VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__inv_8
XTAP_TAPCELL_ROW_11_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_clk_X clkload29/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__mux4_2_A0 hold827/A hold292/A
+ hold470/A hold430/A fanout477/X m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[20\]_sky130_fd_sc_hd__and2_2_X/B
+ sky130_fd_sc_hd__mux4_1
Xm_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold412/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_50_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/A
+ hold644/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__o31a_2_A1_B1 fanout408/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold27/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__and2_2_B fanout436/X hold103/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[2\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold543/X hold1134/A fanout557/X VGND VGND VPWR VPWR hold544/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XFILLER_12_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_71_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout426_X fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload2 clkload2/A VGND VGND VPWR VPWR clkload2/Y sky130_fd_sc_hd__inv_6
XTAP_TAPCELL_ROW_22_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__and2_2
Xm_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold566/X fanout571/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_76_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout408/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold349/A sky130_fd_sc_hd__dfxtp_1
Xfanout250 fanout252/X VGND VGND VPWR VPWR fanout250/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_911 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout261 fanout263/X VGND VGND VPWR VPWR fanout261/X sky130_fd_sc_hd__buf_2
Xfanout272 fanout273/X VGND VGND VPWR VPWR fanout272/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1253/X m_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout602/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout74_X fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout283 fanout283/A VGND VGND VPWR VPWR fanout283/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout294 fanout295/X VGND VGND VPWR VPWR fanout294/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2 m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A2 m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1 m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout473/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout215/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_61_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_matrix\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold128/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[10\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold912/X m_blake2.m_hash256.m_matrix\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout585/X
+ VGND VGND VPWR VPWR hold913/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout300/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold709 hold709/A VGND VGND VPWR VPWR hold709/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout176/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/A1
+ m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/A2 m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/X sky130_fd_sc_hd__o21a_1
XFILLER_48_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A
+ hold653/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold101/X fanout316/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[7\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1045/X m_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout540/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[8\].m_y_buf m_blake2.m_hash256.g_buffer\[8\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[8\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__nand2_2_B fanout433/X hold156/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_A1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_B2
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/X m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X_A1 m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold158/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_56_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__a22o_2_A1 hold260/A fanout294/X
+ fanout405/X hold878/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_19_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__mux2_1_A0 hold352/A m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout383/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__and2_2_B fanout431/X hold174/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_61_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_C1
+ fanout350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X/A1
+ m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X/A2 m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR ANTENNA_13/DIODE sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__and2_2_A/B fanout425/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__o21bai_2_A1 m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__o21bai_2_A1/Y
+ sky130_fd_sc_hd__o21bai_2
XANTENNA_fanout121_A fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout219_A fanout220/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout512/X m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__inv_2
XFILLER_1_918 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A0 hold230/A m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout490_A fanout494/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout235/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1_A
+ fanout301/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__a22o_2_A1 hold366/A fanout187/X
+ fanout195/X hold594/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1041/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/Y m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold69 hold69/A VGND VGND VPWR VPWR hold69/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1 hold823/A fanout382/X
+ fanout186/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__a22o_2_A1 hold467/A fanout191/X
+ fanout200/X hold836/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout256/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[10\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold896/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_S fanout416/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_7_Left_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XFILLER_69_1080 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout182/X m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_4
Xdata\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X data\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata\[2\]_sky130_fd_sc_hd__mux2_1_A1 hold16/X hold15/X fanout598/X VGND VGND VPWR
+ VPWR data\[2\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B fanout498/X hold31/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold226/X m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[11\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[11\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold695/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold541/A fanout53/X fanout81/X m_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_50_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold637/A m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout385/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold1130/A fanout42/X m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_35_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold760/X fanout218/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout245/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1215/A fanout127/X fanout115/X hold931/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1 hold511/A fanout307/X m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/B1
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 VGND VGND VPWR VPWR m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/X
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_63_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_13_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B fanout434/X hold1102/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_15_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_matrix\[14\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1130/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_B m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold517 hold517/A VGND VGND VPWR VPWR hold517/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1262/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_2
Xhold506 hold506/A VGND VGND VPWR VPWR hold506/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X
+ hold416/A fanout352/X fanout183/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__a21o_1
Xhold528 hold528/A VGND VGND VPWR VPWR hold528/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold539 hold539/A VGND VGND VPWR VPWR hold539/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout551/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[13\]\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B fanout206/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_4
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout184/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
Xhold1206 hold1206/A VGND VGND VPWR VPWR hold1206/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1217 hold1217/A VGND VGND VPWR VPWR hold1217/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1239 hold1239/A VGND VGND VPWR VPWR hold1239/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1228 hold1228/A VGND VGND VPWR VPWR hold1228/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hash\[0\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_A fanout402/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ hold427/X fanout216/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_966 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y
+ m_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout88/X
+ fanout116/X hold803/A m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/A3
+ sky130_fd_sc_hd__a221oi_1
Xm_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1098/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__a221o_2_A1_B2 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout336_A fanout341/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__and3_2_A hold307/A fanout465/X fanout376/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XFILLER_55_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold644/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold357/X m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hash\[4\]_sky130_fd_sc_hd__mux2_1_A0_S fanout485/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_60_clk clkload2/A VGND VGND VPWR VPWR clkbuf_leaf_60_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_21_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout420/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__a21o_2_B1/X m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout124_X fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_73_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N/Y
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X hold502/X fanout409/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B fanout493/X m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__xor2_2_B hold979/A hold596/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
XFILLER_0_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout426/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold468/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_40_1404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_C1
+ fanout350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A0 hold62/A m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout513/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold1009/A fanout137/X m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_17_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/B2 hold1004/X fanout588/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold800/X m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_data\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_51_clk clkload3/A VGND VGND VPWR VPWR clkload26/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold342/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold77/A m_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout507/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[22\]_sky130_fd_sc_hd__or2_2_A hold1240/A fanout247/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[22\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_56_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B/Y
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ sky130_fd_sc_hd__a21oi_2
XFILLER_49_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XFILLER_10_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_56_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout289/X m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_52_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout193/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[15\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold549/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__mux2_1_A0 hold776/X m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold922/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1083 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold382/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold859/X m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout156/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_62_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N_sky130_fd_sc_hd__and3_2_X
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/A m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B
+ m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/A_N
+ sky130_fd_sc_hd__and3_1
XFILLER_56_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__or2_2_A hold447/A fanout372/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_42_clk clkload5/A VGND VGND VPWR VPWR clkbuf_leaf_42_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold413/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout232/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X m_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold68/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__xor2_2_B hold617/A hold380/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xhold303 hold303/A VGND VGND VPWR VPWR hold303/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X
+ hold512/A fanout275/X m_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__o21ba_2_A1/X
+ fanout237/X fanout270/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X/B1
+ sky130_fd_sc_hd__a221o_1
Xhold314 hold314/A VGND VGND VPWR VPWR hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 hold325/A VGND VGND VPWR VPWR hold325/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 hold347/A VGND VGND VPWR VPWR hold347/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 hold336/A VGND VGND VPWR VPWR hold336/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold369 hold369/A VGND VGND VPWR VPWR hold369/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2/X
+ sky130_fd_sc_hd__a41o_2
Xm_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold479/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold358 hold358/A VGND VGND VPWR VPWR hold358/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_buffer\[29\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 hold1014/A VGND VGND VPWR VPWR hold1014/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1003 hold1003/A VGND VGND VPWR VPWR hold1003/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1058 hold1058/A VGND VGND VPWR VPWR hold1058/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 hold1047/A VGND VGND VPWR VPWR hold1047/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 hold1036/A VGND VGND VPWR VPWR hold1036/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
Xhold1025 hold1025/A VGND VGND VPWR VPWR hold1025/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout286_A fanout287/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1069 hold1069/A VGND VGND VPWR VPWR hold1069/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_54_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A0 hold55/A m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout519/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout40/X
+ fanout76/X m_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout620_A fanout621/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[57\]_sky130_fd_sc_hd__a21oi_2_A1 hold159/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/X fanout421/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[57\]_sky130_fd_sc_hd__o21a_2_A1/B1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold284/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_33_clk clkload4/A VGND VGND VPWR VPWR clkbuf_leaf_33_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/D m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_652 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3b_2_A_N
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/B1
+ sky130_fd_sc_hd__nand3b_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[6\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout170/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold870 hold870/A VGND VGND VPWR VPWR hold870/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 hold881/A VGND VGND VPWR VPWR hold881/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2
+ fanout293/X m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ fanout356/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2/Y
+ sky130_fd_sc_hd__a211oi_1
Xm_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold967/A fanout86/X fanout98/X hold1209/A m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold892 hold892/A VGND VGND VPWR VPWR hold892/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X hold486/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[12\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1 fanout462/X m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/X
+ sky130_fd_sc_hd__o31a_1
Xm_blake2.m_hash256.m_matrix\[8\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold995/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold880/A fanout32/X fanout76/X m_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout350/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__a21oi_2_B1 fanout446/X m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C/B
+ m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C/C VGND VGND VPWR VPWR
+ m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__a21oi_2_B1/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_input14_A uio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_24_clk clkload1/A VGND VGND VPWR VPWR clkload18/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_matrix\[3\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold698/X hold863/A fanout601/X VGND VGND VPWR VPWR hold699/A sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_45_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y
+ fanout283/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout156/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout283/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ fanout328/X m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B fanout488/X m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_1281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ fanout456/X fanout152/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout482/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA_m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout178/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[2\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_799 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_15_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold1200/A fanout110/X fanout130/X m_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_23_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__xor2_2_A hold1247/A hold438/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A hold270/A m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout283/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold100 hold100/A VGND VGND VPWR VPWR hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout201_A fanout204/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1097/A fanout43/X fanout79/X m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xhold133 hold133/A VGND VGND VPWR VPWR hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A VGND VGND VPWR VPWR hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold122 hold122/A VGND VGND VPWR VPWR hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 hold111/A VGND VGND VPWR VPWR hold111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold177/A VGND VGND VPWR VPWR hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold155/A VGND VGND VPWR VPWR hold155/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold166 hold166/A VGND VGND VPWR VPWR hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout613 fanout614/X VGND VGND VPWR VPWR fanout613/X sky130_fd_sc_hd__buf_2
Xfanout602 fanout603/X VGND VGND VPWR VPWR fanout602/X sky130_fd_sc_hd__buf_2
Xhold199 hold199/A VGND VGND VPWR VPWR hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[1\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold435/X hold378/X fanout557/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold188 hold188/A VGND VGND VPWR VPWR hold188/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold265/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input6_A ui_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/C
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold56/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout289_X fanout289/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold203/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold443/X fanout326/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.ll_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold1235/X fanout167/X m_io.m_config.ll_q\[28\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__a22o_2_A1 hold377/A fanout293/X
+ fanout281/X hold676/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A1
+ fanout487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout284/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__a31o_2_B1_A3
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.g_buffer\[1\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold807/A fanout275/X fanout176/X m_blake2.m_hash256.v_q\[14\]\[31\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout272/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_1107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold276/X
+ fanout165/X m_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X VGND
+ VGND VPWR VPWR hold277/A sky130_fd_sc_hd__o211a_1
XFILLER_46_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X
+ hold1211/A fanout114/X fanout98/X hold1120/A m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y/B
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2/B1
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o2111a_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__xnor2_2_B hold1030/A hold533/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_34_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__mux2_1_A0 hold34/A m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout203/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A/B
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__o21a_2_A1 hold1013/A fanout387/X
+ fanout251/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_47_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout507/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_75_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_47_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__xnor2_2_A hold492/A hold835/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold513/X m_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout543/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[19\]_sky130_fd_sc_hd__or2_2_A hold1105/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[19\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold90/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
Xm_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout161/X m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout611/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_4_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_4_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold183/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout403/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout249_A fanout249/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X
+ hold915/A fanout376/X fanout237/X m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X/A1 sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__and2_2_B fanout436/X hold53/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__and2_2_B_A fanout431/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1082/A fanout91/X fanout150/X m_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__xnor2_2_A hold254/A hold686/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1155/X m_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout550/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout416_A fanout416/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_30_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout204_X fanout204/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[14\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold530/X hold948/A fanout598/X VGND VGND VPWR VPWR hold531/A sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold233/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A0 hold63/A m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout523/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ fanout413/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold331/X hold630/X fanout603/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout421 fanout422/X VGND VGND VPWR VPWR fanout421/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1 hold1190/A fanout275/X
+ fanout176/X m_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__or2_2_A/X fanout270/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xfanout432 fanout434/X VGND VGND VPWR VPWR fanout432/X sky130_fd_sc_hd__buf_2
Xfanout410 fanout412/A VGND VGND VPWR VPWR fanout410/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold971/A sky130_fd_sc_hd__dfxtp_1
Xfanout465 fanout465/A VGND VGND VPWR VPWR fanout465/X sky130_fd_sc_hd__buf_2
Xfanout454 hold409/A VGND VGND VPWR VPWR fanout454/X sky130_fd_sc_hd__buf_2
XFILLER_47_806 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout443 fanout443/A VGND VGND VPWR VPWR fanout443/X sky130_fd_sc_hd__buf_4
Xfanout498 fanout499/X VGND VGND VPWR VPWR fanout498/X sky130_fd_sc_hd__buf_2
Xfanout487 fanout489/X VGND VGND VPWR VPWR fanout487/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__xnor2_2_A hold320/A hold308/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout18/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout476 fanout477/X VGND VGND VPWR VPWR fanout476/X sky130_fd_sc_hd__buf_2
XFILLER_8_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout52/X fanout68/X
+ hold934/A m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_76_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/A1
+ sky130_fd_sc_hd__or4_1
XFILLER_64_89 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/A
+ hold442/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout197/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout83 fanout83/A VGND VGND VPWR VPWR fanout83/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[14\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xfanout50 fanout51/A VGND VGND VPWR VPWR fanout50/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__xor2_2_B hold365/A hold282/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xfanout61 fanout63/X VGND VGND VPWR VPWR fanout61/X sky130_fd_sc_hd__buf_2
Xfanout72 fanout75/A VGND VGND VPWR VPWR fanout72/X sky130_fd_sc_hd__clkbuf_4
Xfanout94 fanout95/A VGND VGND VPWR VPWR fanout94/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout279/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__o21ai_2_A1/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__xnor2_2_A hold1237/A hold997/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1102/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout411/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_36_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold249/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/A1
+ sky130_fd_sc_hd__inv_2
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhash\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A hash\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[7\]_sky130_fd_sc_hd__and2_2_B/B sky130_fd_sc_hd__dfxtp_4
XFILLER_80_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and3_2_C fanout447/X fanout480/X
+ hold64/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XFILLER_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout480/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout196/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1122/X
+ fanout552/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_0_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_53_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1215/A fanout606/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xclkload20 clkload20/A VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__inv_12
Xclkload31 clkload31/A VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__inv_8
Xm_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X/B1
+ m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_11_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A0 hold74/A m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__xnor2_2_A hold550/A hold869/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X hold951/A fanout174/X
+ m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2 hold477/A m_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[28\].m_c_buf/A sky130_fd_sc_hd__a221o_1
XFILLER_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout199_A fanout200/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_1
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR fanout27/A sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold747/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31oi_2_Y
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/A m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X/B
+ m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__a31oi_2
XFILLER_29_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_A fanout371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_820 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout154_X fanout154/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__nand3_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_X fanout419/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload3 clkload3/A VGND VGND VPWR VPWR clkload3/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_22_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X
+ fanout131/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_22_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold890/A fanout112/X fanout120/X m_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_76_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y
+ fanout71/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__o211a_2_A1_A1 m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold1156/A fanout80/X fanout64/X hold1040/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfanout240 fanout240/A VGND VGND VPWR VPWR fanout240/X sky130_fd_sc_hd__buf_4
Xfanout262 fanout263/X VGND VGND VPWR VPWR fanout262/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ fanout452/X fanout454/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_2
Xfanout273 fanout273/A VGND VGND VPWR VPWR fanout273/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__xor2_2_B hold1100/A hold431/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_1
Xfanout251 fanout252/X VGND VGND VPWR VPWR fanout251/X sky130_fd_sc_hd__buf_4
Xfanout284 fanout285/X VGND VGND VPWR VPWR fanout284/X sky130_fd_sc_hd__buf_4
XFILLER_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout295 fanout295/A VGND VGND VPWR VPWR fanout295/X sky130_fd_sc_hd__clkbuf_4
XFILLER_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1060/A fanout59/X fanout71/X hold1007/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_65_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__a211oi_2_A1_A2 fanout283/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout247/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__nor2_4
XFILLER_2_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold331/A fanout147/X fanout123/X m_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold310/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X
+ m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout101/X m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ sky130_fd_sc_hd__o22a_4
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold1167/A fanout146/X fanout122/X m_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D
+ m_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_1326 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__a21oi_2_A1 hold436/A fanout279/X
+ m_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__a22o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__a21oi_2_A1/Y sky130_fd_sc_hd__a21oi_1
XFILLER_80_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout448/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_B2
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_A1
+ fanout266/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X
+ hold1119/A fanout124/X fanout128/X hold702/A m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold733/X VGND VGND VPWR VPWR hold732/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold228/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1135/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold742/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout114_A fanout115/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout345/X m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__a22o_2_A1/X fanout177/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_71_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold230/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout188/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[7\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/B fanout227/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XFILLER_27_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout483_A fanout484/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_69_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_5_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__nor2_2_B fanout490/X hold99/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold806/X m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A hold1159/X
+ VGND VGND VPWR VPWR hold1158/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout271_X fanout271/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_3_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1148/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__mux2_1_A0_A0 m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__and2_2_B fanout442/X hold206/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_73_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A1_S fanout412/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold266/A m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__or2_2_B/X fanout371/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2/A1 fanout227/X VGND VGND VPWR
+ VPWR m_blake2.m_hash256.v_q\[12\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__a22o_2_A1_B2 fanout520/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__or2_2_A hold323/A fanout378/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_8_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout269/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ hold815/X VGND VGND VPWR VPWR hold814/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold172/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2/Y
+ m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__a211oi_2_A1/Y m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout402/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold470/X m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout234/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold775/X fanout223/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A hold365/A m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold314/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold571/X hold563/X fanout589/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold734/X m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout413/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout345/X m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X fanout255/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout194/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold637/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X fanout615/X
+ m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X/B VGND VGND
+ VPWR VPWR m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ hold945/X VGND VGND VPWR VPWR hold944/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_67_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XFILLER_35_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold520/A fanout111/X fanout131/X hold983/A m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__mux2_1_A0 hold235/X hold683/A
+ fanout578/X VGND VGND VPWR VPWR hold236/A sky130_fd_sc_hd__mux2_1
XFILLER_34_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout523/X m_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_63_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__or2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_63_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__a22o_2_A1 hold169/X fanout329/X
+ m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__nand2_2_A hold963/A fanout352/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y
+ fanout194/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout273/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold271/X m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout230/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold384/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__a211o_2_A1_C1 fanout399/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout260/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold680/X hold585/X fanout576/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold507 hold507/A VGND VGND VPWR VPWR hold507/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/A m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/B
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ba_1
Xhold518 hold518/A VGND VGND VPWR VPWR hold518/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold529 hold529/A VGND VGND VPWR VPWR hold529/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_B fanout103/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1080/X m_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout572/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/D
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.g_buffer\[1\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_2
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
XFILLER_48_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1207 hold1207/A VGND VGND VPWR VPWR hold1207/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__o21ai_2_A1 hold1245/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout423/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[14\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold387/X m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout210/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ hold362/X VGND VGND VPWR VPWR hold361/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1218 hold1218/A VGND VGND VPWR VPWR hold1218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_923 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1229 hold1270/A VGND VGND VPWR VPWR hold1229/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold718/X hold873/A fanout574/X VGND VGND VPWR VPWR hold719/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold626/A fanout44/X fanout72/X m_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_hash\[0\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_B m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold404/A m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout395/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout425/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1134 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__a221o_2_A1_A2 m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_C1
+ fanout346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout231_A fanout232/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout329_A fanout330/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1112/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold486/X m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout557/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__mux2_1_A1_A0
+ fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_Y
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_S fanout301/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__a22o_2_A1/X sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__a22o_2_B2 m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ fanout262/X fanout306/X hold276/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A hold194/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold112/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout486_X fanout486/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X/A1
+ fanout343/X VGND VGND VPWR VPWR fanout307/A sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/A
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/Y
+ sky130_fd_sc_hd__nor3_1
XANTENNA_m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold62/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2 m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ fanout264/X fanout307/X hold797/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_45_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold350/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__and2_2_A m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1005/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_40_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold77/X fanout316/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold870/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold631/A fanout147/X fanout151/X m_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout223/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/B sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_55_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold814/A fanout61/X fanout39/X hold898/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout449/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2 m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A1
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 fanout240/X hold1143/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/C1
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/X sky130_fd_sc_hd__o221a_1
Xm_blake2.m_hash256.m_matrix\[5\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold768/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1087/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_7_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B/A
+ VGND VGND VPWR VPWR fanout83/A sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold918/X fanout548/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A hold770/A hold971/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout520/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[11\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold621/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__mux2_1_A1_S fanout214/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__mux2_1_A0 hold61/A m_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_255 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_X m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_S fanout416/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold304 hold304/A VGND VGND VPWR VPWR hold304/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold326 hold326/A VGND VGND VPWR VPWR hold326/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 hold315/A VGND VGND VPWR VPWR hold315/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 hold348/A VGND VGND VPWR VPWR hold348/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold359 hold359/A VGND VGND VPWR VPWR hold359/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 hold337/A VGND VGND VPWR VPWR hold337/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__or2_2_A hold213/A fanout241/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_5_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1004 hold1004/A VGND VGND VPWR VPWR hold1004/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_5_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 hold1015/A VGND VGND VPWR VPWR hold1015/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1048 hold1048/A VGND VGND VPWR VPWR hold1048/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1037 hold1037/A VGND VGND VPWR VPWR hold1037/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 hold1026/A VGND VGND VPWR VPWR hold1026/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 hold1059/A VGND VGND VPWR VPWR hold1059/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout181_A fanout184/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout279_A fanout283/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_22_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold55/X fanout326/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout446_A fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__nor3b_2_Y
+ fanout466/X fanout474/X fanout470/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ sky130_fd_sc_hd__nor3b_4
XFILLER_53_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1211/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[13\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1099/X hold1082/X fanout598/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout613_A fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout234_X fanout234/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_664 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout176/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout401_X fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A/B
+ fanout358/X fanout261/X m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__and3_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold860 hold860/A VGND VGND VPWR VPWR hold860/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 hold882/A VGND VGND VPWR VPWR hold882/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X m_io.m_config.ll_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1064/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2/A1
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
Xhold871 hold871/A VGND VGND VPWR VPWR hold871/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 hold893/A VGND VGND VPWR VPWR hold893/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_10_Left_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout505/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_77_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_904 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold326/X m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ fanout230/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A0 hold178/A m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout504/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold1270/A fanout136/X m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_17_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_c_buf\[14\]_sky130_fd_sc_hd__o22a_2_X hold1035/A fanout175/X
+ m_blake2.m_hash256.g_c_buf\[14\]_sky130_fd_sc_hd__o22a_2_X/B1 fanout253/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[14\].m_c_buf/A sky130_fd_sc_hd__o22a_1
XFILLER_41_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout303/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_45_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold465/X m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout419/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_2
XFILLER_4_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_848 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold845/X fanout551/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0_S fanout299/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold975/A fanout56/X fanout72/X hold946/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_973 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1_A2
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold843/A sky130_fd_sc_hd__dfxtp_1
Xhold101 hold101/A VGND VGND VPWR VPWR hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A VGND VGND VPWR VPWR hold112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold134/A VGND VGND VPWR VPWR hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y/B sky130_fd_sc_hd__a21oi_1
Xhold123 hold123/A VGND VGND VPWR VPWR hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 hold145/A VGND VGND VPWR VPWR hold145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_1360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold167 hold167/A VGND VGND VPWR VPWR hold167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 hold156/A VGND VGND VPWR VPWR hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout603 fanout607/X VGND VGND VPWR VPWR fanout603/X sky130_fd_sc_hd__clkbuf_4
Xfanout614 fanout615/X VGND VGND VPWR VPWR fanout614/X sky130_fd_sc_hd__buf_2
Xhold189 hold189/A VGND VGND VPWR VPWR hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold178 hold178/A VGND VGND VPWR VPWR hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1/X
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1/A1
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A0 hold148/A m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout511/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X
+ hold638/A fanout115/X fanout147/X m_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a221o_1
Xm_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B fanout405/X
+ m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_28_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold514/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout184_X fanout184/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_S fanout222/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2
+ m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B/X
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__a31oi_4
Xm_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_27_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_962 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__or3_2_B fanout407/X hold463/A
+ fanout366/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__or3_2_B/X
+ sky130_fd_sc_hd__or3_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_S fanout232/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0 hold660/X m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_40_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__nor2_2_B_A fanout492/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_1 fanout453/X fanout457/X
+ fanout461/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_1/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_6_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__and3_2_A hold214/A fanout464/X fanout383/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_matrix\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1193/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold968/A fanout140/X fanout120/X data\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
XFILLER_29_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold690 hold690/A VGND VGND VPWR VPWR hold690/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold437/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y fanout270/X m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/X
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XFILLER_79_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold720/A fanout60/X fanout80/X m_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_47_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__nand2_2_B fanout429/X hold225/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold948/X m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout596/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XFILLER_13_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2
+ fanout455/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__or2_2_B fanout488/X hold24/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__xnor2_2_B hold689/A hold588/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_23_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_A_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/D
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B/A
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold957/A fanout56/X fanout44/X hold1066/A m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__xnor2_2_A hold413/A hold575/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_io.cmd\[5\]_sky130_fd_sc_hd__and2b_2_B m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR m_io.cmd\[5\]_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
XANTENNA_m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout144_A fanout147/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_S fanout158/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_S fanout302/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout409_A fanout410/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold100/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold63/X fanout329/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xfanout422 fanout422/A VGND VGND VPWR VPWR fanout422/X sky130_fd_sc_hd__buf_2
XANTENNA_fanout399_X fanout399/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout411 fanout412/X VGND VGND VPWR VPWR fanout411/X sky130_fd_sc_hd__buf_4
Xfanout400 fanout400/A VGND VGND VPWR VPWR fanout400/X sky130_fd_sc_hd__buf_6
Xfanout455 fanout456/X VGND VGND VPWR VPWR fanout455/X sky130_fd_sc_hd__buf_2
Xfanout466 fanout468/A VGND VGND VPWR VPWR fanout466/X sky130_fd_sc_hd__buf_4
Xfanout444 fanout445/A VGND VGND VPWR VPWR fanout444/X sky130_fd_sc_hd__buf_2
Xfanout433 fanout434/X VGND VGND VPWR VPWR fanout433/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout499 fanout500/X VGND VGND VPWR VPWR fanout499/X sky130_fd_sc_hd__clkbuf_4
Xfanout488 fanout489/X VGND VGND VPWR VPWR fanout488/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__a21o_2_X_A1
+ fanout284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout477 fanout477/A VGND VGND VPWR VPWR fanout477/X sky130_fd_sc_hd__buf_4
XFILLER_46_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1/Y
+ sky130_fd_sc_hd__a31oi_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X_sky130_fd_sc_hd__a31o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1/X
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1_sky130_fd_sc_hd__nand2b_2_Y_A_N
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout40 fanout43/A VGND VGND VPWR VPWR fanout40/X sky130_fd_sc_hd__buf_4
XFILLER_30_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.round_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ fanout459/X fanout152/X m_blake2.m_hash256.round_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout482/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xfanout51 fanout51/A VGND VGND VPWR VPWR fanout51/X sky130_fd_sc_hd__clkbuf_2
Xfanout62 fanout63/X VGND VGND VPWR VPWR fanout62/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xfanout73 fanout75/A VGND VGND VPWR VPWR fanout73/X sky130_fd_sc_hd__clkbuf_2
XFILLER_23_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[1\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold397/X hold725/X fanout605/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout95 fanout95/A VGND VGND VPWR VPWR fanout95/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/C
+ sky130_fd_sc_hd__a21o_1
XFILLER_31_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout84 fanout87/A VGND VGND VPWR VPWR fanout84/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_1 hold272/A m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout396/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold619/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold201/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__mux2_1_A0 hold19/A m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout512/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1/C1
+ sky130_fd_sc_hd__clkinv_2
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1032/A fanout58/X fanout54/X m_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_49_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[8\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold950/X m_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout565/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/A
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA_m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout19/X m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[18\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XFILLER_21_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_60_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__and3_2_C_A fanout448/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout416/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout403/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold434/X fanout162/X m_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xclkload10 clkload10/A VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinv_8
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload32 clkload32/A VGND VGND VPWR VPWR clkload32/Y sky130_fd_sc_hd__clkinv_2
Xclkload21 clkload21/A VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__inv_16
Xm_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold71/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_11_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold74/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1133/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XFILLER_68_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold505/X
+ fanout164/X m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__or2_2_A/X fanout617/X VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__o31a_2_A1_A2 fanout385/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A/B sky130_fd_sc_hd__nor2_1
XFILLER_3_1154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout359_A fanout361/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2 m_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout408/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[27\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_34_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and4_2_X
+ fanout449/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/B sky130_fd_sc_hd__and4_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout526_A fanout538/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A0 hold1189/A m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout532/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xclkload4 clkload4/A VGND VGND VPWR VPWR clkload4/X sky130_fd_sc_hd__clkbuf_8
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold1030/X m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_22_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout314_X fanout314/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__a22o_2_A1 hold623/A fanout190/X
+ fanout198/X hold555/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout241 fanout243/X VGND VGND VPWR VPWR fanout241/X sky130_fd_sc_hd__buf_2
Xfanout230 fanout232/A VGND VGND VPWR VPWR fanout230/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_B
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A/C
+ sky130_fd_sc_hd__and2_1
Xfanout274 fanout274/A VGND VGND VPWR VPWR fanout274/X sky130_fd_sc_hd__buf_6
Xfanout263 fanout264/X VGND VGND VPWR VPWR fanout263/X sky130_fd_sc_hd__clkbuf_2
Xfanout252 fanout252/A VGND VGND VPWR VPWR fanout252/X sky130_fd_sc_hd__buf_4
XFILLER_43_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/C
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_31_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__a22o_2_A1 hold446/A fanout188/X
+ fanout196/X hold567/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout296 fanout299/A VGND VGND VPWR VPWR fanout296/X sky130_fd_sc_hd__buf_4
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout178/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout285 fanout288/A VGND VGND VPWR VPWR fanout285/X sky130_fd_sc_hd__buf_4
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout161/X m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout611/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout154/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold1016/A fanout72/X m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_65_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__or2_2_A hold687/A fanout393/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_42_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_61_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X data\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold199/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout419/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__and2_2_A m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_61_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[11\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1063/X m_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout566/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold946/X hold933/X fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xdata\[7\]_sky130_fd_sc_hd__mux2_1_A1 hold300/X hold239/X fanout573/X VGND VGND VPWR
+ VPWR data\[7\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1166/A sky130_fd_sc_hd__dfxtp_1
Xm_io.cmd\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.cmd\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__a32o_2_B2/A2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold916/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold1221/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XFILLER_66_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X
+ fanout468/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X/A3
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X/B1
+ fanout401/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/C
+ sky130_fd_sc_hd__a32o_1
XANTENNA_m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_A1
+ fanout279/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_1299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1207/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout62/X
+ fanout78/X hold1067/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1/A2 m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y/A2
+ fanout427/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1 m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_B2 m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold737/X fanout208/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold769/X m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout301/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout107_A fanout107/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_71_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold512/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__xnor2_2_B hold1185/A hold676/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[12\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold708/X m_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout604/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout16/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout476_A fanout477/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[30\]_sky130_fd_sc_hd__or2_2_A hold196/A fanout247/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[30\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_3_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold688/X m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout126/X
+ fanout94/X m_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B_A
+ fanout288/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[9\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1119/X m_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout564/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout431_X fanout431/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold648/A fanout60/X fanout40/X hold1065/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_78_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__xor2_2_A hold788/A hold753/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A hold1126/X
+ VGND VGND VPWR VPWR hold1223/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold820/X m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout597/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold604/X m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout160/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__a32o_2_A1 hold694/A fanout346/X
+ fanout250/X fanout171/X m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__a32o_2_A1/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_48_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout416/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2
+ fanout287/X m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout280/X fanout359/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold578/X m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_220 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[13\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold861/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A hold312/X
+ VGND VGND VPWR VPWR hold311/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_968 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold965/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A1_S fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_448 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold231/A m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout530/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_63_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout422/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/B fanout227/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold293/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1048 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__or2_2_A hold1247/A fanout362/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold486/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_13_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[10\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold456/X m_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout545/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[15\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ data\[1\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
Xhold508 hold508/A VGND VGND VPWR VPWR hold508/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold519 hold519/A VGND VGND VPWR VPWR hold519/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B hold1255/A
+ hold830/A m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/X
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_29_Left_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold721/X m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout153/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold525/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[2\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold920/A sky130_fd_sc_hd__dfxtp_1
Xhold1219 hold1219/A VGND VGND VPWR VPWR hold1219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_935 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1208 hold1208/A VGND VGND VPWR VPWR hold1208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold404/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
XFILLER_19_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout198/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2
+ m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout501/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold793/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[4\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[4\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1081/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout224_A fanout224/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__a21o_2_A1 hold76/X fanout315/X
+ m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A_1 m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ fanout459/X fanout461/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A_1/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.v_q\[8\]\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold682/X fanout224/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold237/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_48_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_A1
+ fanout285/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_B2
+ fanout279/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold648/X data\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout543/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_matrix\[15\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__mux2_1
Xhash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/X
+ hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout309/X VGND VGND VPWR VPWR hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[3\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout357/X m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__a22o_2_A1/X fanout179/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XFILLER_38_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__or2_2_B fanout487/X hold91/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N/X
+ fanout362/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2/Y
+ sky130_fd_sc_hd__o211ai_1
Xm_blake2.m_hash256.m_matrix\[8\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ hold848/X VGND VGND VPWR VPWR hold1067/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_A
+ m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1 fanout454/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold81/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_S fanout218/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold141/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload2_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_B m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1/B1 sky130_fd_sc_hd__and2b_1
XFILLER_21_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold61/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__o2bb2a_2_A1_N m_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout306/X fanout394/X hold831/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_1_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_18_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/X m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/A2_N
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[14\]\[22\]_sky130_fd_sc_hd__or2_2_A hold387/A fanout383/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[22\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_11_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[0\]_sky130_fd_sc_hd__a211o_2_X_A1 m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[20\].m_c_buf m_blake2.m_hash256.g_buffer\[20\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[20\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xhold316 hold316/A VGND VGND VPWR VPWR hold316/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold814/A fanout121/X fanout148/X m_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1086/X m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout156/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold305 hold305/A VGND VGND VPWR VPWR hold305/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 hold349/A VGND VGND VPWR VPWR hold349/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold338 hold338/A VGND VGND VPWR VPWR hold338/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold327 hold327/A VGND VGND VPWR VPWR hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__o22a_2_A2/B1
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_5_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ hold286/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold1005 hold1005/A VGND VGND VPWR VPWR hold1005/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1016 hold1016/A VGND VGND VPWR VPWR hold1016/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 hold1049/A VGND VGND VPWR VPWR hold1049/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 hold1038/A VGND VGND VPWR VPWR hold1038/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1027 hold1027/A VGND VGND VPWR VPWR hold1027/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B fanout486/X hold97/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_61_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__or2_2_B fanout488/X hold149/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A0 hold921/A m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__xnor2_2_A hold352/A hold717/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout174_A fanout174/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout541/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout341_A fanout342/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N/X
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout439_A fanout441/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdata_v_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X data_v_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout608/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_676 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout292/X m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ fanout356/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout286/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout284/X m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B/X fanout346/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold97/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X hold909/A fanout17/X m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[15\].m_y_buf/A sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xhold861 hold861/A VGND VGND VPWR VPWR hold861/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold850 hold850/A VGND VGND VPWR VPWR hold850/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 hold872/A VGND VGND VPWR VPWR hold872/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1038/X hold1015/X fanout579/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout87_A fanout87/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold883 hold883/A VGND VGND VPWR VPWR hold883/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 hold894/A VGND VGND VPWR VPWR hold894/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__a22o_2_A1 hold392/A fanout290/X
+ fanout278/X hold735/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold190/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_C
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ hold818/X VGND VGND VPWR VPWR hold817/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[27\]_sky130_fd_sc_hd__or2_2_A hold243/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[27\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold483/X hold976/A fanout601/X VGND VGND VPWR VPWR hold484/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold178/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_28_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B fanout489/X hold280/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout42_X fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_c_buf\[11\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A/Y
+ fanout253/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[11\]_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_73_1001 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout295/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_buffer\[6\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_58_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold434/A sky130_fd_sc_hd__dfxtp_1
Xdata\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold199/X fanout308/A VGND VGND VPWR VPWR data\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold566/X m_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout571/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A0 hold237/A m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__xnor2_2_A hold637/A hold834/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__xor2_2_X_X
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_A
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X
+ fanout466/X fanout469/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X/A
+ sky130_fd_sc_hd__and2_1
XFILLER_24_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_1_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout295/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xhold135 hold135/A VGND VGND VPWR VPWR hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold124/A VGND VGND VPWR VPWR hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 hold102/A VGND VGND VPWR VPWR hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A VGND VGND VPWR VPWR hold113/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold157 hold157/A VGND VGND VPWR VPWR hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A VGND VGND VPWR VPWR hold168/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold146 hold146/A VGND VGND VPWR VPWR hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout615 input2/X VGND VGND VPWR VPWR fanout615/X sky130_fd_sc_hd__clkbuf_2
Xfanout604 fanout605/X VGND VGND VPWR VPWR fanout604/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[14\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold179 hold179/A VGND VGND VPWR VPWR hold179/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold148/X fanout323/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__a22o_2_A1_A1 m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_A fanout295/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__nand2_2_B_A fanout437/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout177_X fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold658/A fanout30/X fanout38/X hold1183/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_6_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X
+ m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout100/X m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B/A
+ sky130_fd_sc_hd__o22a_4
XFILLER_27_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout359/X m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__a22o_2_A1/X fanout179/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_54_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold376/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_buffer\[21\].m_y_buf m_blake2.m_hash256.g_buffer\[21\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[21\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_clkbuf_leaf_69_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout289/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.g_buffer\[12\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_6_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_A1 hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[22\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_B
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A0 hold54/A m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold680 hold680/A VGND VGND VPWR VPWR hold680/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold691 hold691/A VGND VGND VPWR VPWR hold691/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1052/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
XFILLER_49_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__xnor2_2_B hold477/A hold504/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__a21o_2_A1_A2 fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1088 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_2
XFILLER_75_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_47_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[3\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold975/X hold957/X fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A hold234/A m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_41_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B
+ fanout444/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_A1/Y VGND
+ VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_51_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_2
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1117/A fanout30/X fanout38/X hold1248/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_4_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout87/X fanout90/X
+ m_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_67_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2_B1 fanout307/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ hold381/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 fanout240/X hold1105/A
+ m_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XFILLER_48_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold735/X m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout413/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_1_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__or2_2_A hold418/A fanout379/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout137_A fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold522/X m_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout604/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload23/A m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout480/A sky130_fd_sc_hd__dfxtp_4
Xm_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__or2_2_A hold389/A fanout373/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout304_A fanout307/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[8\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold702/X hold1049/X fanout562/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold944/A fanout70/X m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xfanout423 fanout424/X VGND VGND VPWR VPWR fanout423/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout401 fanout403/X VGND VGND VPWR VPWR fanout401/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/A
+ hold562/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout412 fanout412/A VGND VGND VPWR VPWR fanout412/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X
+ hold1048/A fanout381/X fanout240/X m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__inv_2_A/Y
+ fanout271/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__o221a_1
Xfanout456 fanout456/A VGND VGND VPWR VPWR fanout456/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout182/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout445 fanout445/A VGND VGND VPWR VPWR fanout445/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout434 fanout443/X VGND VGND VPWR VPWR fanout434/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout294_X fanout294/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout489 fanout500/A VGND VGND VPWR VPWR fanout489/X sky130_fd_sc_hd__buf_4
Xfanout478 fanout480/A VGND VGND VPWR VPWR fanout478/X sky130_fd_sc_hd__clkbuf_4
Xm_io.data_v_early_sky130_fd_sc_hd__and3_2_C hold1/A hold5/A data_v_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.data_v_early_sky130_fd_sc_hd__and3_2_C/X sky130_fd_sc_hd__and3_1
Xfanout467 fanout468/A VGND VGND VPWR VPWR fanout467/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout221/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xblock_first_sky130_fd_sc_hd__a22o_2_B2 fanout485/X block_last_sky130_fd_sc_hd__a22o_2_B2/A2
+ block_last_sky130_fd_sc_hd__a22o_2_B2/B1 hold13/X VGND VGND VPWR VPWR block_first_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_1375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.fsm_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout610/X fanout482/X m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and3_1
Xm_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__or2_2_A hold511/A fanout248/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_14_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout189/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout30 fanout31/A VGND VGND VPWR VPWR fanout30/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1037 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout74 fanout75/A VGND VGND VPWR VPWR fanout74/X sky130_fd_sc_hd__clkbuf_4
Xfanout63 fanout63/A VGND VGND VPWR VPWR fanout63/X sky130_fd_sc_hd__buf_2
XFILLER_11_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout52 fanout55/A VGND VGND VPWR VPWR fanout52/X sky130_fd_sc_hd__clkbuf_4
Xfanout41 fanout43/A VGND VGND VPWR VPWR fanout41/X sky130_fd_sc_hd__buf_2
XFILLER_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout419/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout85 fanout87/A VGND VGND VPWR VPWR fanout85/X sky130_fd_sc_hd__clkbuf_2
Xfanout96 fanout99/A VGND VGND VPWR VPWR fanout96/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold174/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_36_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B
+ fanout476/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold645/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_S fanout221/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_1448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_896 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B fanout489/X m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout188/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_61_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__o22a_2_A1 hold825/A m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ fanout173/X fanout254/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__o22a_1
XANTENNA_data\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1241/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__or2_2_A hold717/A fanout383/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xclkload33 clkload33/A VGND VGND VPWR VPWR clkload33/Y sky130_fd_sc_hd__inv_8
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload22 clkload22/A VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__inv_4
Xclkload11 clkload11/A VGND VGND VPWR VPWR clkload11/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[13\]\[2\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold724/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2
+ fanout266/X m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout400/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_68_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/X m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2/A2_N
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_1
XFILLER_60_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__o31a_2_A1_A3 fanout249/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_852 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold151/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_844 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1197/X fanout604/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout135/X
+ fanout123/X m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A_A m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold1189/X fanout330/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout421_A fanout422/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__o21a_2_X
+ hold961/A fanout381/X fanout185/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__o21a_1
Xclkload5 clkload5/A VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_6
XANTENNA_fanout519_A fanout524/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout307_X fanout307/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1011/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[14\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1065/X m_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout543/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_796 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_S fanout228/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__a22o_2_A1 hold678/A fanout292/X
+ fanout286/X hold596/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold714/A sky130_fd_sc_hd__dfxtp_1
Xfanout231 fanout232/A VGND VGND VPWR VPWR fanout231/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A_A m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout473/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout220 fanout220/A VGND VGND VPWR VPWR fanout220/X sky130_fd_sc_hd__buf_4
Xfanout242 fanout243/X VGND VGND VPWR VPWR fanout242/X sky130_fd_sc_hd__clkbuf_2
Xfanout264 fanout265/X VGND VGND VPWR VPWR fanout264/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout253 fanout254/X VGND VGND VPWR VPWR fanout253/X sky130_fd_sc_hd__buf_4
Xfanout297 fanout299/A VGND VGND VPWR VPWR fanout297/X sky130_fd_sc_hd__buf_2
Xfanout275 fanout276/A VGND VGND VPWR VPWR fanout275/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold107/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_47_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout286 fanout287/X VGND VGND VPWR VPWR fanout286/X sky130_fd_sc_hd__clkbuf_4
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold540/X VGND VGND VPWR VPWR hold539/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold476/A m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout386/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_A_N
+ m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout360/X m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X fanout257/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold35/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A0 hold474/A m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout512/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold572/A fanout275/X m_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout185/X fanout271/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout35/X fanout71/X
+ hold821/A m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XFILLER_24_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold689/X m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_61_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__nand2_2_A hold1018/A fanout343/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold702/A fanout77/X fanout72/X hold943/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_S fanout303/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X
+ fanout269/X m_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__and4_1
Xm_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold496/X m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2_B1_sky130_fd_sc_hd__nand2_2_Y
+ fanout463/X fanout373/X VGND VGND VPWR VPWR fanout240/A sky130_fd_sc_hd__nand2_2
Xm_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y/B
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ hold516/A m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D
+ m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__a22o_2_A1 hold545/A fanout190/X
+ fanout198/X hold1069/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xblock_first_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__inv_2_Y block_last_sky130_fd_sc_hd__a32o_2_B2/A1
+ VGND VGND VPWR VPWR block_first_sky130_fd_sc_hd__a32o_2_B2/A1 sky130_fd_sc_hd__clkinv_2
Xm_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2 m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ fanout262/X fanout307/X hold360/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ sky130_fd_sc_hd__a22oi_1
Xm_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__nand2_2_A hold1226/A fanout343/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ hold622/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2/A1
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold299/X m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout230/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold260/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_72_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_72_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A2 m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.g_buffer\[6\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[14\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold308/X m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout212/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[12\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold708/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ fanout462/X fanout152/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout482/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold979/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold399/A m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout367/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout540/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_69_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold838/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/A fanout219/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y
+ fanout168/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR fanout71/A sky130_fd_sc_hd__nor2_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_21_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout371_A fanout399/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_S fanout214/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold61/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_72_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold366/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C_C
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1186/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_37_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout257_X fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout41/X
+ fanout76/X m_blake2.m_hash256.m_matrix\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_63_clk clkload2/A VGND VGND VPWR VPWR clkload23/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout415/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.m_matrix\[1\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold826/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold826/A fanout25/X m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_78_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold467/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.v_q\[13\]\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold285/X fanout207/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold867/A fanout61/X fanout41/X hold1071/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__a221o_2_B2_C1 fanout268/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1214/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
XFILLER_3_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold1002/A fanout132/X fanout121/X data\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout17/X m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[30\].m_y_buf/A sky130_fd_sc_hd__o32a_1
Xm_io.m_config.ll_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold307/X fanout164/X m_io.m_config.ll_q\[24\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold485/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold795/X fanout220/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout72_X fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold78/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[3\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[3\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1032/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold888/A sky130_fd_sc_hd__dfxtp_1
XFILLER_43_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_67_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__a32o_2_B1/A2
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold231/X fanout335/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold1157/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_54_clk clkload3/A VGND VGND VPWR VPWR clkload27/A sky130_fd_sc_hd__clkbuf_8
XFILLER_15_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout241/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_63_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold528/X
+ fanout161/X m_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X VGND
+ VGND VPWR VPWR hold529/A sky130_fd_sc_hd__o211a_1
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1243/A fanout577/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/A2
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X fanout406/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_16_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR hold1224/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout349/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold471/X m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold509 hold509/A VGND VGND VPWR VPWR hold509/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[5\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A hold1184/X
+ VGND VGND VPWR VPWR hold1183/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__xnor2_2_A hold779/A m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_buffer\[14\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N/X
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A0 hold278/A m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout536/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold421/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A0 hold252/A m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout519/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1209 hold1209/A VGND VGND VPWR VPWR hold1209/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__or2_2_A hold908/A fanout364/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold807/X m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_S fanout203/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold172/A m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_45_clk clkload3/A VGND VGND VPWR VPWR clkload25/A sky130_fd_sc_hd__clkbuf_8
XFILLER_34_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__a32o_2_B1/A3
+ sky130_fd_sc_hd__nand2_1
XFILLER_34_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1
+ fanout284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A fanout166/X m_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout619/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_S fanout419/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold722/A fanout51/X fanout47/X hold811/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_A fanout218/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A data\[7\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold300/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[9\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold938/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold1013/X m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout155/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/B2
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__and2_2_A hold1008/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
XFILLER_56_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1 m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_77_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_36_clk clkload4/A VGND VGND VPWR VPWR clkload33/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__xor2_2_B hold388/A hold436/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
XFILLER_77_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold1017/A m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__or2_2_B/X fanout395/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1079/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2_A1
+ hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_B1
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout90/X
+ fanout114/X hold1248/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_1318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1066/X fanout547/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold817/A fanout124/X fanout88/X hold771/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X
+ hold457/A fanout383/X fanout176/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/A
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X_A2 m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A0 hold197/A m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout529/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold513/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_S fanout221/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clkload1/A VGND VGND VPWR VPWR clkload19/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A_Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout181/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold754/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold889/X m_blake2.m_hash256.m_matrix\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout565/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_18_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ sky130_fd_sc_hd__and2b_1
XFILLER_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1_A1_N
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1215/X hold1213/X fanout606/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR fanout236/A sky130_fd_sc_hd__nor2_2
Xm_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A/B
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A/C
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/X VGND
+ VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_matrix\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold974/X hold931/X fanout601/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold564/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__or2_2_B fanout493/X hold63/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xhold306 hold306/A VGND VGND VPWR VPWR hold306/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold317 hold317/A VGND VGND VPWR VPWR hold317/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR fanout107/A sky130_fd_sc_hd__and4_2
Xhold328 hold328/A VGND VGND VPWR VPWR hold328/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 hold339/A VGND VGND VPWR VPWR hold339/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_buffer\[24\].m_c_buf m_blake2.m_hash256.g_buffer\[24\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[24\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold574/A fanout88/X fanout120/X m_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X
+ fanout190/X m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o2bb2a_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__a21oi_2_A1/B1 sky130_fd_sc_hd__and2_1
Xhold1006 hold1006/A VGND VGND VPWR VPWR hold1006/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1017 hold1017/A VGND VGND VPWR VPWR hold1017/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hash\[4\]_sky130_fd_sc_hd__mux2_1_A0_A0 hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1039 hold1039/A VGND VGND VPWR VPWR hold1039/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1028 hold1028/A VGND VGND VPWR VPWR hold1028/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold921/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout604/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__o41a_2_B1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ fanout451/X fanout456/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B/D
+ sky130_fd_sc_hd__o41a_1
XANTENNA_fanout167_A fanout168/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_18_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_35_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A_B m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_983 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[7\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold923/X hold889/X fanout567/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout334_A fanout335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold1007/A fanout111/X fanout115/X hold1177/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/X fanout610/X input6/X VGND VGND VPWR VPWR m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_B
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/A3
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_B/X
+ sky130_fd_sc_hd__or3_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold1051/A fanout48/X m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/A2
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_66_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold862 hold862/A VGND VGND VPWR VPWR hold862/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 hold851/A VGND VGND VPWR VPWR hold851/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 hold873/A VGND VGND VPWR VPWR hold873/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold840 hold840/A VGND VGND VPWR VPWR hold840/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xhold884 hold884/A VGND VGND VPWR VPWR hold884/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 hold895/A VGND VGND VPWR VPWR hold895/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X
+ hold668/A fanout87/X m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X/A
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout229/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_48_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout295/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0 hold535/X m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout299/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold45/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout157/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ hold884/X VGND VGND VPWR VPWR hold883/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout303/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold566/A fanout109/X fanout141/X hold826/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_hash\[3\]_sky130_fd_sc_hd__mux2_1_A0_X hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X
+ hold802/A fanout101/X m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A1 sky130_fd_sc_hd__o22a_2
XFILLER_16_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__a221o_2_A1 hold800/A fanout276/X
+ fanout176/A m_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__or2_2_A/X fanout272/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_57_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold680/A fanout125/X m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_58_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__or2_2_B_A fanout487/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1140/A fanout34/X fanout78/X m_blake2.m_hash256.m_matrix\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__or2_2_A hold759/A fanout175/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_80_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold237/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B
+ fanout344/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ fanout276/A sky130_fd_sc_hd__and3_2
XPHY_EDGE_ROW_66_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B
+ m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_23_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_706 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__or2_2_B fanout495/X hold67/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_75_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__xnor2_2_A hold271/A hold526/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_A m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold103 hold103/A VGND VGND VPWR VPWR hold103/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hash_v_sky130_fd_sc_hd__a211o_2_X_C1 fanout478/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold125 hold125/A VGND VGND VPWR VPWR hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A VGND VGND VPWR VPWR hold114/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout425/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold306/A sky130_fd_sc_hd__dfxtp_1
Xhold158 hold158/A VGND VGND VPWR VPWR hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkload8/A sky130_fd_sc_hd__clkbuf_8
Xhold147 hold147/A VGND VGND VPWR VPWR hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 hold136/A VGND VGND VPWR VPWR hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 hold169/A VGND VGND VPWR VPWR hold169/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout605 fanout606/X VGND VGND VPWR VPWR fanout605/X sky130_fd_sc_hd__clkbuf_4
Xfanout616 fanout621/X VGND VGND VPWR VPWR fanout616/X sky130_fd_sc_hd__buf_2
XFILLER_59_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__o21bai_2_A2
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__o21bai_4
Xm_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__xnor2_2_A hold404/A hold372/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout284_A fanout285/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
XFILLER_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_A1
+ fanout418/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__a21o_2_B1/X m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A/B
+ sky130_fd_sc_hd__and2_1
XFILLER_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold871/X hold803/X fanout546/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__and3_2_A hold204/A fanout464/X fanout395/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__inv_2_A hold1237/A VGND VGND VPWR
+ VPWR m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__clkinv_2
XFILLER_23_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout415/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold377/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_40_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_buffer\[25\].m_y_buf m_blake2.m_hash256.g_buffer\[25\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[25\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold274/A sky130_fd_sc_hd__dfxtp_1
Xm_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__mux2_1_X
+ m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q input15/X fanout1/A VGND VGND VPWR VPWR
+ m_io.cmd\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X/B sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold661/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_2_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__a221o_2_A1 hold429/A m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ m_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__or2_2_A/X fanout171/X m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__o21a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[16\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold670 hold670/A VGND VGND VPWR VPWR hold670/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold54/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_9_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold681 hold681/A VGND VGND VPWR VPWR hold681/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold692 hold692/A VGND VGND VPWR VPWR hold692/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1057/A fanout134/X fanout122/X hold752/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_65_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1212/X m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input12_A uio_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/B
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A_X fanout412/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_47_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout98/X fanout150/X
+ hold621/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_26_791 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_c_buf\[4\]_sky130_fd_sc_hd__a211o_2_X hold971/A fanout174/A
+ m_blake2.m_hash256.g_c_buf\[4\]_sky130_fd_sc_hd__a211o_2_X/B1 m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__a32o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[4\].m_c_buf/A sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__mux2_1_A0 hold23/A m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout534/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__and2_2_B fanout428/X hold54/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_12_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_B_sky130_fd_sc_hd__a311o_2_X
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A2
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C/B
+ sky130_fd_sc_hd__a311o_1
Xm_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A0 hold182/A m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold897/X hold826/X fanout571/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout141/X
+ fanout93/X m_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout49/X fanout53/X
+ m_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__and3_2_B ANTENNA_11/DIODE
+ m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_1
XFILLER_58_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[3\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout541/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1259/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_Q
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_A fanout500/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__or2_2_A hold753/A fanout392/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xfanout413 fanout414/X VGND VGND VPWR VPWR fanout413/X sky130_fd_sc_hd__buf_4
XFILLER_28_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout402 fanout403/X VGND VGND VPWR VPWR fanout402/X sky130_fd_sc_hd__clkbuf_4
Xfanout446 fanout448/X VGND VGND VPWR VPWR fanout446/X sky130_fd_sc_hd__buf_4
XANTENNA_input4_A ui_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout424 fanout427/X VGND VGND VPWR VPWR fanout424/X sky130_fd_sc_hd__clkbuf_2
Xfanout457 fanout458/A VGND VGND VPWR VPWR fanout457/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout435 fanout443/X VGND VGND VPWR VPWR fanout435/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout479 fanout480/A VGND VGND VPWR VPWR fanout479/X sky130_fd_sc_hd__clkbuf_2
Xfanout468 fanout468/A VGND VGND VPWR VPWR fanout468/X sky130_fd_sc_hd__buf_2
XANTENNA_fanout287_X fanout287/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_76_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X hash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6/D sky130_fd_sc_hd__a21o_1
XFILLER_70_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout621_X fanout621/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout31 fanout31/A VGND VGND VPWR VPWR fanout31/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout20 fanout23/X VGND VGND VPWR VPWR fanout20/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold784/A fanout124/X fanout97/X m_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout42 fanout43/A VGND VGND VPWR VPWR fanout42/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_42_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout64 fanout67/A VGND VGND VPWR VPWR fanout64/X sky130_fd_sc_hd__buf_4
Xfanout53 fanout55/A VGND VGND VPWR VPWR fanout53/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout75 fanout75/A VGND VGND VPWR VPWR fanout75/X sky130_fd_sc_hd__clkbuf_2
Xfanout86 fanout87/A VGND VGND VPWR VPWR fanout86/X sky130_fd_sc_hd__clkbuf_4
Xfanout97 fanout99/A VGND VGND VPWR VPWR fanout97/X sky130_fd_sc_hd__clkbuf_2
XFILLER_13_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__a2bb2o_2_A1_N/B2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ sky130_fd_sc_hd__or3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ data\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout61/X m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XFILLER_49_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold736/X fanout572/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1/B
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_801 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B fanout424/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XFILLER_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__a22o_2_A1/B1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__o21bai_2_A1/Y m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/X
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3_2_B
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3_2_B/A
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3_2_B/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B fanout499/X hold203/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xclkload34 clkload34/A VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__inv_6
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload12 clkload12/A VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__clkinvlp_4
XTAP_TAPCELL_ROW_11_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload23 clkload23/A VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__inv_16
XFILLER_55_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_53_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_68_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold287/X m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_Y m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout247_A fanout248/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout414_A fanout416/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload6 clkload6/A VGND VGND VPWR VPWR clkload6/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_76_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout202_X fanout202/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1 hold489/A fanout295/X
+ m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__a22o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1/X
+ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_76_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y
+ hash\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0 m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__nand2_1
XFILLER_69_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold321/X m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout210 fanout211/X VGND VGND VPWR VPWR fanout210/X sky130_fd_sc_hd__buf_4
Xfanout232 fanout232/A VGND VGND VPWR VPWR fanout232/X sky130_fd_sc_hd__clkbuf_4
Xfanout221 fanout222/X VGND VGND VPWR VPWR fanout221/X sky130_fd_sc_hd__buf_4
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout477/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold832/A sky130_fd_sc_hd__dfxtp_1
Xfanout243 fanout248/A VGND VGND VPWR VPWR fanout243/X sky130_fd_sc_hd__clkbuf_2
Xfanout265 fanout265/A VGND VGND VPWR VPWR fanout265/X sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_31_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y/B sky130_fd_sc_hd__nand2b_1
Xm_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__xnor2_2_A hold743/A hold330/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xfanout254 fanout254/A VGND VGND VPWR VPWR fanout254/X sky130_fd_sc_hd__clkbuf_8
XFILLER_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout276 fanout276/A VGND VGND VPWR VPWR fanout276/X sky130_fd_sc_hd__buf_2
Xfanout298 fanout299/X VGND VGND VPWR VPWR fanout298/X sky130_fd_sc_hd__buf_4
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout287 fanout288/X VGND VGND VPWR VPWR fanout287/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_A1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout62_A fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout170/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold476/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_4_0_clk_X clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1175/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X
+ m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold76/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold619/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold665/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold517/X m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout158/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_65_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold474/X fanout317/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1202/A fanout542/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/B sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_753 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold193/A fanout142/X fanout95/X hold445/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2
+ fanout266/A m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout400/A fanout389/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ sky130_fd_sc_hd__o221a_1
Xm_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1 hold502/A fanout402/X
+ m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__a22o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_13_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold803/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1163/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[4\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold686/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold272/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[0\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold508/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout596/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_1443 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold325/A m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout372/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__o21bai_2_A1/Y m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/X
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y/B
+ sky130_fd_sc_hd__a21o_1
XFILLER_34_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold519/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout235/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2
+ fanout190/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout181/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.m_matrix\[2\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[2\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold641/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout534/X m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold420/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold666/X m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1056/A fanout110/X fanout150/X hold1256/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X
+ m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold399/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_A2 fanout100/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold42/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__mux2_1_A1_A1 m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout197_A fanout200/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__a22o_2_A1 hold550/A fanout192/X
+ fanout200/X hold627/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR fanout59/A sky130_fd_sc_hd__nor2_2
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[6\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold346/X m_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout570/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold165/X fanout327/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold324/X m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout531_A fanout538/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkload23/A m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__o21a_2_X
+ hold822/A fanout369/X fanout176/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.v_q\[8\]\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold837/X fanout221/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_78_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout417_X fanout417/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout157/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold454/A m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout397/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[30\]_sky130_fd_sc_hd__or2_2_A hold383/A fanout392/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[30\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1136/A fanout128/X fanout96/X m_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1071/X m_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout563/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_16_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_26_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_13_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold649/X fanout604/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[13\]\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold869/X fanout206/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout279/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold169/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold93/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold278/X fanout340/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold189/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__mux2_1_A1_S fanout228/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold252/X fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_1455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold161/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold855/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[3\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[3\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1000/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_B2
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/C m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1 m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_53_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold172/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold755/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout190/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A1
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A2
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A3
+ fanout100/X m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o32ai_4
XANTENNA_m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout184/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A1_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__or2_2_A hold797/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__and2_2_B fanout436/X hold412/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[5\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold736/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold418/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or4_2_A/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout112_A fanout115/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload23/A m_blake2.m_hash256.g_buffer\[20\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold276/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B_A fanout497/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold361/X hold493/A fanout548/X VGND VGND VPWR VPWR hold362/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ fanout457/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A0 hold106/A m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout504/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout417/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout579_A fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_block_data.data_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__mux2_1_X
+ fanout308/X block_last_sky130_fd_sc_hd__a32o_2_B2/A3 hold5/A VGND VGND VPWR VPWR
+ m_io.m_block_data.data_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B_A fanout434/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold936/A fanout138/X m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout255/X m_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout380/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR fanout212/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout25_A fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__a22o_2_A1/B1 sky130_fd_sc_hd__xnor2_1
XFILLER_21_892 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout255/X m_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout367/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold369/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
XFILLER_4_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__nand2_2_Y
+ fanout610/X m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/A2 VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold197/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[29\]_sky130_fd_sc_hd__o22a_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1 hold1262/A fanout357/X
+ fanout262/X m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold259/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout273/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout64/X
+ fanout36/X hold768/A m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_hash\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__and3_2_B_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold307 hold307/A VGND VGND VPWR VPWR hold307/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__a211o_2_A1 hold767/A fanout282/X
+ m_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__a22o_2_A1/X fanout386/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold329 hold329/A VGND VGND VPWR VPWR hold329/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold318 hold318/A VGND VGND VPWR VPWR hold318/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2
+ fanout295/X m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B/X fanout350/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2/Y
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout155/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A0 hold144/A m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X/A1
+ hash_v_sky130_fd_sc_hd__a211o_2_X/A2 hold185/A fanout606/X VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[28\].m_c_buf m_blake2.m_hash256.g_buffer\[28\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[28\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xhold1018 hold1018/A VGND VGND VPWR VPWR hold1018/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold536/A fanout87/X fanout119/X hold1036/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xhold1007 hold1007/A VGND VGND VPWR VPWR hold1007/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 hold1029/A VGND VGND VPWR VPWR hold1029/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1146/X fanout543/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold196/X fanout167/X m_io.m_config.ll_q\[22\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_39_756 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1/B
+ fanout249/X VGND VGND VPWR VPWR fanout194/A sky130_fd_sc_hd__nor2_2
XFILLER_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A ANTENNA_8/DIODE m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_22_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout327_A fanout330/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold905/A sky130_fd_sc_hd__dfxtp_1
Xhold830 hold830/A VGND VGND VPWR VPWR hold830/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X
+ hold369/A fanout126/X fanout134/X m_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a221o_1
Xhold863 hold863/A VGND VGND VPWR VPWR hold863/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold841 hold841/A VGND VGND VPWR VPWR hold841/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold852 hold852/A VGND VGND VPWR VPWR hold852/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold874 hold874/A VGND VGND VPWR VPWR hold874/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__nor2_2_A_A fanout465/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold885 hold885/A VGND VGND VPWR VPWR hold885/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 hold896/A VGND VGND VPWR VPWR hold896/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout484_X fanout484/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B_A fanout489/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1055/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout181/X m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_51_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_S fanout201/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X
+ m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1/B
+ VGND VGND VPWR VPWR fanout55/A sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold630/A fanout54/X fanout34/X hold841/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ fanout252/X m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[11\]\[31\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout172/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_28_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__nand2b_2_B/Y m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__xnor2_2_A hold343/A hold724/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_49_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.g_buffer\[17\].m_y_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_13_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold224/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__a31o_2_A3 fanout446/X fanout479/X
+ hold107/A fanout512/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_45_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout28_X fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout406/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A0 hold227/A m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold620/X fanout576/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold201/X fanout166/X m_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_58_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__xnor2_2_A hold604/A hold547/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1006/A fanout60/X fanout73/X m_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y fanout177/X m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__a21oi_2
Xm_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__xnor2_2_B hold1142/A hold734/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__a211o_2_A1 hold570/A fanout282/X
+ m_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__a22o_2_A1/X fanout387/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_23_1403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__nor2_2_A fanout465/A fanout344/X
+ VGND VGND VPWR VPWR fanout265/A sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B_B m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_A0
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B_A m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2_A1
+ hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1138/X m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout154/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold127/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2_B2 m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y fanout273/X m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_30_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold115 hold115/A VGND VGND VPWR VPWR hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold1108/A fanout84/X fanout88/X m_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xhold126 hold126/A VGND VGND VPWR VPWR hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold104 hold104/A VGND VGND VPWR VPWR hold104/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A_B m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold159 hold159/A VGND VGND VPWR VPWR hold159/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1
+ fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold148 hold148/A VGND VGND VPWR VPWR hold148/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__xnor2_2_A hold721/A hold556/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold137 hold137/A VGND VGND VPWR VPWR hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout606 fanout607/X VGND VGND VPWR VPWR fanout606/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold150/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
Xfanout617 fanout621/X VGND VGND VPWR VPWR fanout617/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_clkload14_A clkload14/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_339 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_S fanout224/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1167/X fanout594/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout277_A fanout278/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_1_A1
+ fanout413/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1084/X fanout570/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_14_Left_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout232_X fanout232/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1053 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1031 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B fanout486/X hold810/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_68_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold563/X m_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout601/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_2_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_buffer\[29\].m_y_buf m_blake2.m_hash256.g_buffer\[29\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[29\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xhold660 hold660/A VGND VGND VPWR VPWR hold660/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1066/A fanout136/X fanout140/X hold1202/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_9_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold671 hold671/A VGND VGND VPWR VPWR hold671/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A
+ fanout487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold693 hold693/A VGND VGND VPWR VPWR hold693/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold682 hold682/A VGND VGND VPWR VPWR hold682/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[0\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold894/X hold1162/A fanout550/X VGND VGND VPWR VPWR hold895/A sky130_fd_sc_hd__mux2_1
XFILLER_79_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1 m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/X
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2/B1
+ m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_715 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_47_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XFILLER_33_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold386/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A hold1160/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
XFILLER_13_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout195/X m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout187/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A_A m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold488/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout596/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xdata\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold12/X fanout308/X VGND VGND VPWR VPWR data\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_S fanout228/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold182/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_A2_sky130_fd_sc_hd__and2_2_X_X
+ fanout174/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1_C1
+ fanout178/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/A
+ sky130_fd_sc_hd__inv_2
XFILLER_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A/C
+ sky130_fd_sc_hd__nand2_1
XFILLER_23_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold932/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X hold1100/A m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[25\].m_c_buf/A sky130_fd_sc_hd__a22o_1
XFILLER_17_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[7\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A/B fanout206/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout521/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__xor2_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout302/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A0 hold31/A m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1 m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout307/X m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1/B1 m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B_A fanout434/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_30_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[5\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1085/X m_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout564/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__o21a_2_A1 hold763/A fanout386/X
+ fanout253/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xfanout414 fanout416/A VGND VGND VPWR VPWR fanout414/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_28_1133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout403 fanout406/A VGND VGND VPWR VPWR fanout403/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__or2_2_B_A fanout485/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout447 fanout448/X VGND VGND VPWR VPWR fanout447/X sky130_fd_sc_hd__buf_4
Xfanout425 fanout427/X VGND VGND VPWR VPWR fanout425/X sky130_fd_sc_hd__clkbuf_2
Xfanout436 fanout443/X VGND VGND VPWR VPWR fanout436/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__nand2_2_A_B m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout458 fanout458/A VGND VGND VPWR VPWR fanout458/X sky130_fd_sc_hd__clkbuf_2
Xfanout469 fanout470/X VGND VGND VPWR VPWR fanout469/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1006/X hold886/X fanout576/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout182_X fanout182/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout561_A fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout353/X m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__a22o_2_A1/X fanout178/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__a21o_2_A1_A2 fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout216/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand3_2_C/B
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X/A1
+ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout447_X fanout447/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR fanout19/A sky130_fd_sc_hd__or2_2
XFILLER_15_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout345/X m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__a22o_2_A1/X fanout177/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
Xfanout21 fanout23/X VGND VGND VPWR VPWR fanout21/X sky130_fd_sc_hd__buf_2
XFILLER_80_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout614_X fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout43 fanout43/A VGND VGND VPWR VPWR fanout43/X sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_42_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout54 fanout55/A VGND VGND VPWR VPWR fanout54/X sky130_fd_sc_hd__clkbuf_4
Xfanout65 fanout67/A VGND VGND VPWR VPWR fanout65/X sky130_fd_sc_hd__buf_2
Xfanout32 fanout35/A VGND VGND VPWR VPWR fanout32/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout98 fanout99/A VGND VGND VPWR VPWR fanout98/X sky130_fd_sc_hd__clkbuf_4
Xfanout87 fanout87/A VGND VGND VPWR VPWR fanout87/X sky130_fd_sc_hd__buf_2
XFILLER_10_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout76 fanout79/A VGND VGND VPWR VPWR fanout76/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__a22o_2_A1 hold711/A fanout293/X
+ fanout287/X hold468/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_X clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ hold1068/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold423/A m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout390/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold490 hold490/A VGND VGND VPWR VPWR hold490/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_S fanout214/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__mux2_1_A0 hold18/A m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1190 hold1190/A VGND VGND VPWR VPWR hold1190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__nand2_2_B/Y
+ fanout266/X fanout372/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_72_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
XFILLER_61_857 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_B m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_S fanout415/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold989/A fanout65/X fanout68/X m_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_4
Xclkload13 clkload13/A VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__inv_6
Xclkload24 clkload24/A VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__inv_16
XFILLER_9_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__a22o_2_A1 hold406/A fanout191/X
+ fanout199/X hold922/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1/Y
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N/Y
+ sky130_fd_sc_hd__o21bai_2
XFILLER_79_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold673/X m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0_S
+ fanout520/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold556/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold676/X m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_824 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout188/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout196/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_1359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[11\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1113/X hold989/X fanout548/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload7 clkload7/A VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_fanout407_A fanout408/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[11\]\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold477/X fanout220/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold327/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_76_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_76_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__and2_2_B fanout430/X hold86/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_30_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xena_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__inv_2_Y fanout609/X VGND VGND VPWR
+ VPWR ena_sky130_fd_sc_hd__or2_2_B/A sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout352/X m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__nor2_1
XFILLER_65_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold623/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A0 hold469/A m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout211 fanout212/X VGND VGND VPWR VPWR fanout211/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_A2_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/C m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1/A2
+ sky130_fd_sc_hd__or2_1
Xfanout200 fanout200/A VGND VGND VPWR VPWR fanout200/X sky130_fd_sc_hd__buf_2
Xfanout222 fanout224/A VGND VGND VPWR VPWR fanout222/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold995/A fanout77/X m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_35_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_S fanout201/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout244 fanout248/X VGND VGND VPWR VPWR fanout244/X sky130_fd_sc_hd__clkbuf_2
Xfanout255 fanout258/A VGND VGND VPWR VPWR fanout255/X sky130_fd_sc_hd__buf_4
Xfanout233 fanout234/X VGND VGND VPWR VPWR fanout233/X sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_31_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold391/A sky130_fd_sc_hd__dfxtp_1
Xfanout299 fanout299/A VGND VGND VPWR VPWR fanout299/X sky130_fd_sc_hd__buf_4
Xfanout277 fanout278/X VGND VGND VPWR VPWR fanout277/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout266 fanout266/A VGND VGND VPWR VPWR fanout266/X sky130_fd_sc_hd__buf_6
Xfanout288 fanout288/A VGND VGND VPWR VPWR fanout288/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold223/X m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A/B fanout207/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/A
+ hold1217/A hold652/A VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_2
Xm_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold446/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold480/X m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_S fanout417/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1174/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_1270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold617/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout24/X m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2 fanout531/X hold143/A
+ m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/B1 m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__or2_2_B fanout494/X hold382/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold804/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[12\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold1104/X VGND VGND VPWR VPWR hold1170/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold368/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold341/X m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout418/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_38_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold1149/A fanout58/X fanout46/X hold914/A m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold325/X fanout410/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A_B
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1051/A fanout96/X fanout148/X hold1175/A m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_4_1455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout407/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
XFILLER_33_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold598/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold297/X m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.g_buffer\[19\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold373/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_block_data.data_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_io.m_block_data.data_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold5/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__o21a_2_A1 hold996/A fanout386/X
+ fanout170/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B fanout490/X hold253/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold918/X m_blake2.m_hash256.m_matrix\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout549/X
+ VGND VGND VPWR VPWR hold919/A sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_71_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[12\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1244/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold133/A m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout504/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y fanout270/X m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1120/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_S fanout221/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold256/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_927 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[0\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1233/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_A
+ fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1119/A fanout33/X fanout41/X m_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_Q
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1
+ fanout301/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout357_A fanout361/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout229/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout524_A fanout539/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_78_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout155/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold936/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold298/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold454/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold11/A fanout62/X fanout34/X m_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__a221o_2_A1 hold1019/A fanout275/X
+ m_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__or2_2_A/X fanout185/X fanout270/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2 m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/A1_N
+ m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/A2_N m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout58_X fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A hold1116/X
+ VGND VGND VPWR VPWR hold1115/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_67_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[3\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1015/X hold491/X fanout567/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[8\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1230/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__xor2_2_B hold1021/A hold681/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_52_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[8\]\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold835/X fanout222/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout132/X
+ fanout140/X hold378/A m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A2
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_13_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B_A fanout486/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_67_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_2_Left_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold634/A fanout129/X fanout149/X hold1063/A m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ fanout423/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XFILLER_7_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__mux4_2_A0_S0 fanout477/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[6\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold911/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_matrix\[15\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ VGND VGND VPWR VPWR fanout43/A sky130_fd_sc_hd__nor2_2
XFILLER_48_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload21/A m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1180/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/Y m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_A_N
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1/X m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_A_N/X
+ sky130_fd_sc_hd__and2b_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XFILLER_26_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold653/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/X sky130_fd_sc_hd__xor2_1
XFILLER_74_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout157/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[8\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_blake2.m_hash256.m_matrix\[8\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold790/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_hash\[4\]_sky130_fd_sc_hd__mux2_1_A0_X hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_B2
+ fanout400/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_A1
+ fanout266/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout302/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold938/A fanout126/X fanout94/X m_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A fanout449/X fanout454/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_4
Xm_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold121/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_73_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold180/A sky130_fd_sc_hd__dfxtp_1
Xdata_idx\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X hold1/X VGND VGND VPWR
+ VPWR data_idx\[0\]_sky130_fd_sc_hd__and4_2_B/C sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[8\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold847/X m_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout593/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__and3_2_C_A fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout105_A fanout107/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold173/X fanout330/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold106/X fanout312/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout401/X m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__o22a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__nand2_2_B fanout428/X hold290/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold994/A fanout146/X fanout122/X m_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1146/A fanout108/X fanout132/X hold1050/A m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_72_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold798/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold783/A fanout96/X m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold131/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__o21a_2_A1 m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B/A
+ fanout362/X fanout407/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A0 hold118/A m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__or2_2_A hold276/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_56_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout501/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_43_1033 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_7_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__xnor2_2_A hold476/A hold1035/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_47_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_A2
+ fanout103/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N/Y
+ sky130_fd_sc_hd__o21bai_1
XFILLER_35_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[7\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold923/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold929/X fanout589/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__inv_2_A m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR hash\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__inv_2
XFILLER_71_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold202/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_687 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__o21bai_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold308 hold308/A VGND VGND VPWR VPWR hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ hold1008/X m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout424/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout196/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold136/A sky130_fd_sc_hd__dfxtp_1
Xhold319 hold319/A VGND VGND VPWR VPWR hold319/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[9\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[9\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold750/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ hold4/A m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold144/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold766/A fanout135/X fanout99/X hold929/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1019 hold1019/A VGND VGND VPWR VPWR hold1019/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1008 hold1008/A VGND VGND VPWR VPWR hold1008/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__xnor2_2_A hold299/A hold1083/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout182/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[4\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold943/X hold853/X fanout568/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1206/X m_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout562/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B
+ fanout471/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1/B
+ VGND VGND VPWR VPWR fanout192/A sky130_fd_sc_hd__nor2_4
XFILLER_61_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1095 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_data\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold360/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A0 hold65/A m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout512/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout222_A fanout224/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout549/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ data\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout60/X fanout52/X m_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold820 hold820/A VGND VGND VPWR VPWR hold820/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__xnor2_2_A hold399/A hold1043/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold831 hold831/A VGND VGND VPWR VPWR hold831/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold842 hold842/A VGND VGND VPWR VPWR hold842/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout108_X fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold853 hold853/A VGND VGND VPWR VPWR hold853/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 hold864/A VGND VGND VPWR VPWR hold864/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 hold875/A VGND VGND VPWR VPWR hold875/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 hold886/A VGND VGND VPWR VPWR hold886/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold897 hold897/A VGND VGND VPWR VPWR hold897/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_51_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout477_X fanout477/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__xnor2_2_B hold825/A hold688/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__inv_2_A m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ VGND VGND VPWR VPWR fanout47/A sky130_fd_sc_hd__nor2_2
XFILLER_45_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold16/A fanout62/X fanout70/X hold606/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold392/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_49_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1209/A fanout50/X fanout46/X m_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_49_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold146/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_45_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/X VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/A1_N sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold227/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout299/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B
+ fanout407/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_58_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_801 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout29/X
+ fanout37/X m_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A hold1246/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_1
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_1/Y
+ sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__or2_2_B fanout484/X hold960/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold739/A fanout586/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkload0_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[14\]\[2\]_sky130_fd_sc_hd__mux2_1_A0 hold822/X m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.g_buffer\[23\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
XFILLER_56_1279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[3\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold1154/X VGND VGND VPWR VPWR hold1153/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A0 hold120/A m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hash_v_sky130_fd_sc_hd__a211o_2_X_A1 fanout463/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__xnor2_2_A hold471/A hold978/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2_A2 fanout260/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__a22oi_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_8_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold105 hold105/A VGND VGND VPWR VPWR hold105/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout278/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold116 hold116/A VGND VGND VPWR VPWR hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold127 hold127/A VGND VGND VPWR VPWR hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold149/A VGND VGND VPWR VPWR hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_A1
+ fanout285/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold138 hold138/A VGND VGND VPWR VPWR hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__a22o_2_A1/B1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__or2_1
XFILLER_28_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhash\[4\]_sky130_fd_sc_hd__mux2_1_A0 hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout485/X VGND VGND VPWR VPWR hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_4
Xfanout607 fanout608/X VGND VGND VPWR VPWR fanout607/X sky130_fd_sc_hd__clkbuf_2
Xfanout618 fanout621/X VGND VGND VPWR VPWR fanout618/X sky130_fd_sc_hd__buf_2
XFILLER_28_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout159/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold962/X m_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout540/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout172_A fanout173/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xblock_last_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X fanout610/X block_last_sky130_fd_sc_hd__a32o_2_B2/X
+ VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_A_N_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout437_A fanout442/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout409/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout225_X fanout225/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_40_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__xnor2_2_A hold1013/A hold678/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_9_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold650 hold650/A VGND VGND VPWR VPWR hold650/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 hold672/A VGND VGND VPWR VPWR hold672/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 hold661/A VGND VGND VPWR VPWR hold661/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout289/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold683 hold683/A VGND VGND VPWR VPWR hold683/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold694 hold694/A VGND VGND VPWR VPWR hold694/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout286/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout85_A fanout87/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout176/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2/X
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1/X
+ sky130_fd_sc_hd__a21bo_4
Xm_blake2.m_hash256.g_buffer\[10\].m_c_buf m_blake2.m_hash256.g_buffer\[10\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[10\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout40_X fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold1064/X fanout167/X m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ sky130_fd_sc_hd__o21ai_2
XFILLER_25_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold1192/A fanout26/X m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold959/A fanout28/X m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XFILLER_51_1143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout279/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_2
Xm_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold98/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_68_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__nand2b_2
XFILLER_27_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_19_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__o2bb2a_2_A1_N m_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout304/X fanout370/X hold1194/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_36_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold933/X hold415/X fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold928/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__xnor2_2_B hold795/A hold608/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__xnor2_2_B/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold31/X fanout340/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A2
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A2/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_34_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A2
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_30_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout404 fanout406/X VGND VGND VPWR VPWR fanout404/X sky130_fd_sc_hd__buf_4
Xfanout448 fanout448/A VGND VGND VPWR VPWR fanout448/X sky130_fd_sc_hd__clkbuf_8
Xfanout426 fanout427/X VGND VGND VPWR VPWR fanout426/X sky130_fd_sc_hd__clkbuf_4
Xm_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A fanout162/X m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout616/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__mux2_1_A0 hold401/A m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout369/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xfanout415 fanout416/X VGND VGND VPWR VPWR fanout415/X sky130_fd_sc_hd__buf_4
XFILLER_28_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout437 fanout442/X VGND VGND VPWR VPWR fanout437/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold950/A fanout129/X fanout133/X hold1015/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xfanout459 fanout460/A VGND VGND VPWR VPWR fanout459/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout175_X fanout175/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__mux2_1_A1_S fanout323/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xblock_first_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A block_first_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__o211a_2_A1 m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__o211a_2_A1/X sky130_fd_sc_hd__o211a_1
XANTENNA_fanout342_X fanout342/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout22 fanout23/X VGND VGND VPWR VPWR fanout22/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X
+ m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or3b_2_B/C_N
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout55 fanout55/A VGND VGND VPWR VPWR fanout55/X sky130_fd_sc_hd__buf_2
Xfanout33 fanout35/A VGND VGND VPWR VPWR fanout33/X sky130_fd_sc_hd__clkbuf_2
Xfanout44 fanout47/A VGND VGND VPWR VPWR fanout44/X sky130_fd_sc_hd__clkbuf_4
Xfanout99 fanout99/A VGND VGND VPWR VPWR fanout99/X sky130_fd_sc_hd__clkbuf_2
Xfanout66 fanout67/A VGND VGND VPWR VPWR fanout66/X sky130_fd_sc_hd__clkbuf_4
Xfanout77 fanout79/A VGND VGND VPWR VPWR fanout77/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold1142/X m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xfanout88 fanout91/A VGND VGND VPWR VPWR fanout88/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ hold862/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold335/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__xnor2_2_A hold579/A hold561/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold977/X VGND VGND VPWR VPWR hold976/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold423/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold917/X hold727/X fanout576/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold480 hold480/A VGND VGND VPWR VPWR hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_78_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold491 hold491/A VGND VGND VPWR VPWR hold491/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B_A m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout88_X fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold500/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold448/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A hold657/X
+ VGND VGND VPWR VPWR hold656/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold1180 hold1180/A VGND VGND VPWR VPWR hold1180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1191 hold1191/A VGND VGND VPWR VPWR hold1191/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold533/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1_A
+ fanout407/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout271/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xnor2_1
XFILLER_53_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold984/X hold1081/A fanout569/X VGND VGND VPWR VPWR hold985/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__xor2_2_B hold916/A hold327/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold372/X m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout210/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload14 clkload14/A VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinv_2
Xclkload25 clkload25/A VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinvlp_4
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y/A
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y/B
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y/C
+ VGND VGND VPWR VPWR ANTENNA_3/DIODE sky130_fd_sc_hd__nor3_2
XTAP_TAPCELL_ROW_11_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout198/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1039/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout281/X m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B/X fanout355/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[1\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold976/X m_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout605/X
+ VGND VGND VPWR VPWR hold977/A sky130_fd_sc_hd__mux2_1
XFILLER_47_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold450/A m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout366/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__nor2_2_B fanout490/X hold168/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_buffer\[11\].m_y_buf m_blake2.m_hash256.g_buffer\[11\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[11\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__xnor2_2_Y_B
+ m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_980 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1042 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__or2_2_B fanout490/X hold198/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_58_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1131/X fanout593/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold510/X m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout414/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__a32o_2_B1 fanout534/X m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__a32o_2_B1/A2
+ m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__a32o_2_B1/A3 hold10/X fanout338/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_51_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ sky130_fd_sc_hd__and2b_1
Xclkload8 clkload8/A VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__bufinv_16
XANTENNA_m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B_A fanout486/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XFILLER_30_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold57/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout302_A fanout303/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhash\[4\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B fanout403/X hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hash\[4\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_65_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_B1_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__and2_1
XFILLER_69_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__nand2_2_A hold906/A fanout353/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold469/X fanout327/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold245/X m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout230/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xfanout201 fanout204/X VGND VGND VPWR VPWR fanout201/X sky130_fd_sc_hd__buf_4
Xm_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2 m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ fanout259/X fanout304/X hold434/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ sky130_fd_sc_hd__a22oi_1
Xfanout212 fanout212/A VGND VGND VPWR VPWR fanout212/X sky130_fd_sc_hd__buf_2
Xfanout223 fanout224/X VGND VGND VPWR VPWR fanout223/X sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_2
Xfanout245 fanout246/X VGND VGND VPWR VPWR fanout245/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1213/A fanout127/X fanout147/X hold1076/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout256 fanout258/A VGND VGND VPWR VPWR fanout256/X sky130_fd_sc_hd__buf_2
Xfanout234 fanout236/A VGND VGND VPWR VPWR fanout234/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__xnor2_2
Xfanout278 fanout279/X VGND VGND VPWR VPWR fanout278/X sky130_fd_sc_hd__clkbuf_4
Xfanout267 fanout267/A VGND VGND VPWR VPWR fanout267/X sky130_fd_sc_hd__buf_6
XTAP_TAPCELL_ROW_31_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold678/A sky130_fd_sc_hd__dfxtp_1
Xfanout289 fanout290/X VGND VGND VPWR VPWR fanout289/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_66_clk clkload0/A VGND VGND VPWR VPWR clkbuf_leaf_66_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X hold311/A fanout19/X m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[2\].m_y_buf/A sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_2
XANTENNA_fanout48_A fanout51/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_65_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold828/A m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout384/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__o21a_2_A1 hold1265/A fanout364/X
+ fanout171/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold442/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__and2_2_B fanout439/X hold129/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__o21ai_2_A1/A2 m_blake2.m_hash256.block_idx_plus_one_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A0 hold833/A m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_matrix\[5\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold931/X hold749/X fanout601/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__or2_2_A hold1042/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_65_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__a211o_2_A1 hold533/A fanout281/X
+ m_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__a22o_2_A1/X fanout389/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1_A2_sky130_fd_sc_hd__or2_2_X
+ fanout362/X fanout254/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ sky130_fd_sc_hd__or2_4
XFILLER_19_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[1\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[1\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold397/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold545/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_57_clk clkload3/A VGND VGND VPWR VPWR clkbuf_leaf_57_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_4_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_A
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__a211o_2_A1 hold704/A fanout284/X
+ m_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__a22o_2_A1/X fanout363/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_14_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__mux2_1_A0 hold388/X m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout236/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold972/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_S fanout208/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold729/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold864/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__xnor2_2_A hold555/A hold535/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold751/X m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1002/X hold984/X fanout569/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold133/X fanout312/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_29_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold801/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2/A1
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2/X
+ sky130_fd_sc_hd__o21ba_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_S fanout213/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout18/X m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[8\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XFILLER_25_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput1 ena VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_48_clk clkload4/A VGND VGND VPWR VPWR clkbuf_leaf_48_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout558/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_A1_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/A1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold778/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold302/X m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.g_buffer\[25\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout138_X fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1143/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__a221o_2_A1 hold612/A fanout351/X
+ fanout263/X m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y
+ fanout156/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A0 hold44/A m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_X
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_1406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__nor2_2_Y_B
+ m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_S fanout156/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A0 hold810/A m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout511/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_10_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y
+ fanout274/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold653/X m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout95/A sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_54_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_0_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_39_clk clkload5/A VGND VGND VPWR VPWR clkbuf_leaf_39_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
XFILLER_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold349/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_2_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ hold1205/X VGND VGND VPWR VPWR hold1009/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_1_A1
+ fanout418/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold849/A fanout138/X fanout142/X hold553/A m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__mux4_2_A0_S1 m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_S fanout204/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X block_last_sky130_fd_sc_hd__a22o_2_B2/X
+ VGND VGND VPWR VPWR fanout465/A sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__and2_2_A/B fanout423/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__a22o_2_A1 hold34/X fanout322/X
+ m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__a22o_2_A1/B1 fanout515/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a22o_1
XFILLER_47_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B/B
+ fanout320/X m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold980/A fanout108/X fanout128/X m_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold171/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold575/X fanout223/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR fanout23/A sky130_fd_sc_hd__nor2_1
XFILLER_34_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A0 hold114/A m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout214/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout287/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_4
XTAP_TAPCELL_ROW_73_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__and3_2_C_B fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_66_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2/X
+ fanout379/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2/X
+ sky130_fd_sc_hd__o211a_1
Xm_io.cmd\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X fanout1/X fanout609/X
+ input12/X VGND VGND VPWR VPWR m_io.cmd\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and3_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout300/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_728 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1247/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout255_X fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_62_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout49/X fanout53/X
+ m_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XFILLER_13_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout422_X fanout422/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold66/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__or2_2_B_A fanout494/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold118/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_56_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout508/X m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XFILLER_49_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__mux2_1_A0/X
+ m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B/B fanout318/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_S fanout222/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[14\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1074/X m_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout583/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold651/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1415 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__xor2_2_X
+ fanout466/X fanout471/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__xor2_4
XFILLER_28_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold867/X fanout565/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__xnor2_2_A hold517/A hold987/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_44_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[29\]_sky130_fd_sc_hd__o22a_2_A1_A2 m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_16_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1 fanout461/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/C
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B/X fanout401/X fanout468/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1/X
+ sky130_fd_sc_hd__o311a_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2_B1_sky130_fd_sc_hd__and3b_2_X
+ fanout470/X fanout474/X fanout466/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1
+ sky130_fd_sc_hd__and3b_2
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold309 hold309/A VGND VGND VPWR VPWR hold309/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__xor2_2_A hold594/A hold660/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold957/X hold883/X fanout548/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__and3_2_B hold1161/A
+ m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_2
XFILLER_39_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1009 hold1009/A VGND VGND VPWR VPWR hold1009/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__xnor2_2_A hold325/A hold827/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout55/X fanout67/X
+ m_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_739 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_35_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1083 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1_B1
+ fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold553/A fanout26/X m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A hold216/X VGND VGND VPWR
+ VPWR m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__inv_2_Y
+ fanout463/X VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X/A1
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/D
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold65/X fanout320/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout61/X fanout77/X
+ hold634/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout215_A fanout216/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
Xhold821 hold821/A VGND VGND VPWR VPWR hold821/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold810 hold810/A VGND VGND VPWR VPWR hold810/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[11\]_sky130_fd_sc_hd__nor2_2_A_B fanout377/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xhold843 hold843/A VGND VGND VPWR VPWR hold843/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold854 hold854/A VGND VGND VPWR VPWR hold854/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 hold832/A VGND VGND VPWR VPWR hold832/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 hold865/A VGND VGND VPWR VPWR hold865/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold876 hold876/A VGND VGND VPWR VPWR hold876/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold898 hold898/A VGND VGND VPWR VPWR hold898/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 hold887/A VGND VGND VPWR VPWR hold887/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__a31o_2_B1 hold1160/A
+ m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B
+ m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_51_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__a211o_2_A1 hold504/A fanout288/X
+ m_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__a22o_2_A1/X fanout378/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_4_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__xnor2_2_A hold324/A hold1145/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_66_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold443/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_49_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X/A1
+ fanout175/X m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X/B1 fanout254/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[9\].m_c_buf/A sky130_fd_sc_hd__o22a_1
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_S fanout302/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1 m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout307/X m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1/B1 m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_45_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout283/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold826/X m_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout571/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold614/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A0 hold70/A m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout520/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_58_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1 m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold966/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A3 m_io.cmd\[2\]_sky130_fd_sc_hd__nor2_2_A/Y
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/X VGND VGND VPWR VPWR fanout248/A
+ sky130_fd_sc_hd__and3_2
XANTENNA_m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_S
+ fanout371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__xnor2_2_A hold454/A m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_26_Left_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_19_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__and2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblock_last_sky130_fd_sc_hd__a22o_2_B2_B1_sky130_fd_sc_hd__nor2_2_Y fanout422/A block_last_sky130_fd_sc_hd__a22o_2_B2/A2
+ VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__a22o_2_B2/B1 sky130_fd_sc_hd__nor2_1
XFILLER_23_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[4\]_sky130_fd_sc_hd__a211o_2_X_A2 fanout174/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_35_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold14/A fanout62/X fanout42/X m_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_411 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold154/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_32_967 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold120/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0 hold315/A hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X
+ fanout379/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X/A
+ ANTENNA_6/DIODE VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__or2_1
XFILLER_30_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a221o_2_B1
+ fanout444/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_3/X m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1 m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/A
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold117 hold117/A VGND VGND VPWR VPWR hold117/X sky130_fd_sc_hd__dlygate4sd3_1
Xhash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
XPHY_EDGE_ROW_44_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold106 hold106/A VGND VGND VPWR VPWR hold106/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__a31o_2_A3_B1 fanout520/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold128 hold128/A VGND VGND VPWR VPWR hold128/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 hold139/A VGND VGND VPWR VPWR hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xfanout608 fanout608/A VGND VGND VPWR VPWR fanout608/X sky130_fd_sc_hd__buf_2
XFILLER_63_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout619 fanout620/X VGND VGND VPWR VPWR fanout619/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__a211o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_S fanout213/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold601/X fanout592/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ sky130_fd_sc_hd__nor3_1
Xm_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__xor2_2_A hold548/A hold612/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_B2 fanout173/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_53_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A0 hold91/A m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout513/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[14\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold574/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold772/A fanout140/X fanout92/X hold1039/A m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_S fanout413/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
XFILLER_33_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A0 hold108/A m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout528/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout332_A fanout342/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__a21oi_2_B1/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_2
XANTENNA_m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_62_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout218_X fanout218/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout120_X fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X hold835/A fanout174/X
+ m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1 hold665/A m_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[24\].m_c_buf/A sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A hold590/X
+ VGND VGND VPWR VPWR hold589/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold651 hold651/A VGND VGND VPWR VPWR hold651/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold640 hold640/A VGND VGND VPWR VPWR hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold662 hold662/A VGND VGND VPWR VPWR hold662/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold673 hold673/A VGND VGND VPWR VPWR hold673/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold684 hold684/A VGND VGND VPWR VPWR hold684/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 hold695/A VGND VGND VPWR VPWR hold695/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold896/X fanout567/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout543/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_buffer\[14\].m_c_buf m_blake2.m_hash256.g_buffer\[14\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[14\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/A1
+ fanout16/X m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/B1 m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[5\].m_y_buf/A sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.m_matrix\[4\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold839/X hold624/X fanout602/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_4
XPHY_EDGE_ROW_80_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1/B1 m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nor2_2
XFILLER_51_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X
+ hold781/A fanout98/X m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X/C1
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X/D1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X/B
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__nand2_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1_B2
+ fanout188/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_S fanout201/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_48_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_672 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X
+ fanout269/X m_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__and4_1
XFILLER_64_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout417/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__and2_2_B fanout428/X hold147/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1049/A fanout33/X fanout65/X hold421/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_17_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1009/X hold1204/A fanout568/X VGND VGND VPWR VPWR hold1205/A sky130_fd_sc_hd__mux2_1
XFILLER_20_904 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X
+ m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_30_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/A2
+ sky130_fd_sc_hd__and2_1
XFILLER_67_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold270/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout549/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_2
XFILLER_67_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout405 fanout406/X VGND VGND VPWR VPWR fanout405/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout427 fanout427/A VGND VGND VPWR VPWR fanout427/X sky130_fd_sc_hd__buf_4
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/B1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1122/A fanout80/X fanout44/X hold1134/A m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xfanout438 fanout442/X VGND VGND VPWR VPWR fanout438/X sky130_fd_sc_hd__clkbuf_2
Xfanout416 fanout416/A VGND VGND VPWR VPWR fanout416/X sky130_fd_sc_hd__buf_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout449 fanout449/A VGND VGND VPWR VPWR fanout449/X sky130_fd_sc_hd__buf_2
XFILLER_58_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1172/X fanout540/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y
+ fanout307/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout282_A fanout283/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout168_X fanout168/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold997/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1120/X fanout581/X
+ VGND VGND VPWR VPWR hold1121/A sky130_fd_sc_hd__mux2_1
Xhash\[2\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2 fanout401/X hash\[2\]_sky130_fd_sc_hd__mux2_1_A1/X
+ m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__and2_2_B/X fanout285/X fanout345/X
+ VGND VGND VPWR VPWR hash\[2\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2/Y
+ sky130_fd_sc_hd__a221oi_1
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold513/A fanout48/X fanout68/X hold1045/A m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout256/X m_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout373/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_1155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout23 fanout23/A VGND VGND VPWR VPWR fanout23/X sky130_fd_sc_hd__buf_2
Xfanout34 fanout35/A VGND VGND VPWR VPWR fanout34/X sky130_fd_sc_hd__clkbuf_4
Xfanout56 fanout59/A VGND VGND VPWR VPWR fanout56/X sky130_fd_sc_hd__buf_4
XANTENNA_fanout335_X fanout335/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout45 fanout47/A VGND VGND VPWR VPWR fanout45/X sky130_fd_sc_hd__clkbuf_2
Xfanout67 fanout67/A VGND VGND VPWR VPWR fanout67/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[12\]\[3\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1048/X fanout228/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xfanout78 fanout79/A VGND VGND VPWR VPWR fanout78/X sky130_fd_sc_hd__clkbuf_4
Xfanout89 fanout91/A VGND VGND VPWR VPWR fanout89/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__nand2_2_B fanout432/X hold95/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__o311a_2_A1/X
+ m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X/C
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold687/X m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold851/A sky130_fd_sc_hd__dfxtp_1
XFILLER_46_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_S fanout224/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1175/A fanout64/X fanout36/X hold778/A m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xhold470 hold470/A VGND VGND VPWR VPWR hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 hold481/A VGND VGND VPWR VPWR hold481/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold707/X m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold492 hold492/A VGND VGND VPWR VPWR hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_Q
+ m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold526/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold621/A fanout66/X m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_79_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__a22o_2_A1/B1
+ sky130_fd_sc_hd__xnor2_1
Xhold1170 hold1170/A VGND VGND VPWR VPWR hold1170/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input10_A ui_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1181 hold1181/A VGND VGND VPWR VPWR hold1181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1192 hold1192/A VGND VGND VPWR VPWR hold1192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout229/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__a21oi_2_A1_A2 fanout279/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_848 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1_B
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout385/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__o22a_2_A2 fanout501/X hold147/A
+ m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__o22a_2_A2/B1 m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
Xm_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__or2_2_A/A fanout167/X m_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout618/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_matrix\[15\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[15\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1006/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[12\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1206/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold603/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold527/X m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xclkload15 clkload15/A VGND VGND VPWR VPWR clkload15/X sky130_fd_sc_hd__clkbuf_4
Xm_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y
+ hash\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0 m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__nand2_1
XFILLER_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload26 clkload26/A VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__inv_8
Xm_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/X
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y/C
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold492/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2/X
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold450/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ hold935/X VGND VGND VPWR VPWR hold934/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1/B1 sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B/B
+ fanout321/X m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_buffer\[15\].m_y_buf m_blake2.m_hash256.g_buffer\[15\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[15\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout202/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold588/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold3/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_51_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xnor2_1
XANTENNA_m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2
+ fanout163/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload9 clkload9/A VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__inv_8
XFILLER_20_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold820/A fanout110/X fanout130/X hold1179/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout128_A fanout131/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/D
+ m_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold254/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold355/A m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout390/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout247/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout596/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout213 fanout216/X VGND VGND VPWR VPWR fanout213/X sky130_fd_sc_hd__buf_4
Xfanout202 fanout203/X VGND VGND VPWR VPWR fanout202/X sky130_fd_sc_hd__buf_4
XANTENNA_fanout497_A fanout500/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y_Y
+ fanout266/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout246 fanout247/X VGND VGND VPWR VPWR fanout246/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout224 fanout224/A VGND VGND VPWR VPWR fanout224/X sky130_fd_sc_hd__buf_4
Xfanout235 fanout236/X VGND VGND VPWR VPWR fanout235/X sky130_fd_sc_hd__buf_4
XANTENNA_input2_A rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout268 fanout269/A VGND VGND VPWR VPWR fanout268/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout285_X fanout285/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout257 fanout258/X VGND VGND VPWR VPWR fanout257/X sky130_fd_sc_hd__clkbuf_4
Xfanout279 fanout283/A VGND VGND VPWR VPWR fanout279/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_31_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_31_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[11\]\[23\]_sky130_fd_sc_hd__a211o_2_A1 m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/A
+ fanout172/X m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__a22o_2_B1/X fanout253/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[23\]_sky130_fd_sc_hd__o311a_2_X/B1
+ sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout158/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout352/X m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__a22o_2_A1/X fanout180/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XFILLER_54_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout173/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2/X
+ m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout404/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a22o_2
Xm_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold320/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[2\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1066/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold828/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_21_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold129/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold833/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1071/X
+ fanout563/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_1010 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold951/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B/B
+ fanout317/X m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1237/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__xor2_2_A hold1157/A hold687/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2
+ hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ sky130_fd_sc_hd__a21bo_1
XFILLER_24_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[8\]\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold834/X fanout223/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2
+ fanout274/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_815 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X
+ fanout408/X fanout355/X m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ sky130_fd_sc_hd__and3_4
XFILLER_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1185/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[2\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1066/X hold1050/X fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold763/X fanout223/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold409/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR fanout228/A sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold343/X m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold74/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A0 hold746/A m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout532/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout411/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1 m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_9_1324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput2 rst_n VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_matrix\[9\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1213/X m_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout607/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B
+ fanout304/X m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR fanout186/A sky130_fd_sc_hd__nor2_2
XFILLER_49_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold550/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_1
XFILLER_65_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[21\]_sky130_fd_sc_hd__or2_2_A hold291/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[21\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold113/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XFILLER_40_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold184/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X
+ m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1259/X m_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout569/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__o21a_2_A1 hold872/A fanout378/X
+ fanout173/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[4\]_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout412_A fanout412/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold667/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold44/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B
+ m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y/B m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/X
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__nor3_1
Xm_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold712/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout200_X fanout200/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[9\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1215/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout74/X m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload21/A m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold810/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout101/X hold852/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B/A
+ sky130_fd_sc_hd__o32a_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout141/X
+ fanout117/X m_blake2.m_hash256.m_matrix\[13\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout91/A sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_54_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold909/X hold1233/A fanout577/X VGND VGND VPWR VPWR hold910/A sky130_fd_sc_hd__mux2_1
XFILLER_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold415/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout60_A fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_675 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_A
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_26_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.g_buffer\[31\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_26_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xuio_out_sky130_fd_sc_hd__buf_2_X uio_out_sky130_fd_sc_hd__buf_2_X/A VGND VGND VPWR
+ VPWR uio_out[3] sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
Xm_io.m_config.ll_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_io.m_config.ll_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold986/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A0 hold1022/A m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A_1_Y fanout295/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A0 hold1263/A m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__o21a_2_A1 hold1044/A fanout365/X
+ fanout250/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1_A2_sky130_fd_sc_hd__or2_2_X_X
+ m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_52_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/X
+ m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__xnor2_2_A hold423/A hold901/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_61_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XFILLER_76_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_943 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/A
+ m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/B m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/X sky130_fd_sc_hd__or3_1
XFILLER_34_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout286/X m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout280/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold229/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_77_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[5\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold690/X hold781/A fanout585/X VGND VGND VPWR VPWR hold691/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold114/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2/A1
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_4
XFILLER_31_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout195_A fanout197/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout347/X m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__a22o_2_A1/X fanout177/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold676/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_951 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_B fanout354/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__nor3b_2_Y
+ fanout466/X fanout469/X fanout475/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ sky130_fd_sc_hd__nor3b_4
XFILLER_52_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__and2_2_A/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout150_X fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout248_X fanout248/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout66/X
+ fanout74/X hold958/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_36_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout415_X fanout415/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A0 hold1012/A m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout511/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X
+ fanout147/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[1\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/X
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_56_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y
+ m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.m_matrix\[13\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold803/X hold574/X fanout549/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y_A
+ m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold766/X fanout601/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout63_X fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold1076/A fanout55/X fanout35/X hold1213/A m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ sky130_fd_sc_hd__or2_1
XFILLER_54_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_2
Xm_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_11_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21ba_2_X
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/A m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o21ba_1
XFILLER_7_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout189/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout394/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout196/X m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout188/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.g_buffer\[28\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[14\]\[7\]_sky130_fd_sc_hd__mux2_1_A0 hold1092/X m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout210/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold789/X m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1259/A fanout568/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X
+ m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1204/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__xnor2_2_A hold297/A hold1181/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_17_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[5\]_sky130_fd_sc_hd__mux2_1_A1_A0 hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/X
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[17\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_17_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout537/X m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XFILLER_61_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/B
+ fanout357/X fanout261/X m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ fanout269/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_50_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1223/X
+ fanout565/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__xnor2_2_B hold241/A hold666/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold800 hold800/A VGND VGND VPWR VPWR hold800/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout110_A fanout111/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold811 hold811/A VGND VGND VPWR VPWR hold811/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 hold855/A VGND VGND VPWR VPWR hold855/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 hold822/A VGND VGND VPWR VPWR hold822/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 hold833/A VGND VGND VPWR VPWR hold833/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold844 hold844/A VGND VGND VPWR VPWR hold844/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__xnor2_2_A hold801/A hold595/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold866 hold866/A VGND VGND VPWR VPWR hold866/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1068 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_X
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold877 hold877/A VGND VGND VPWR VPWR hold877/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold888 hold888/A VGND VGND VPWR VPWR hold888/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold899 hold899/A VGND VGND VPWR VPWR hold899/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__a21oi_2_B1_A1 fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout198_X fanout198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X
+ hold376/A fanout374/X fanout193/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/B
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_51_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XFILLER_44_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_28_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__or2_2_B_A fanout485/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__or2_2_A hold1143/A fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_49_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_965 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B/X m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_73_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/A
+ hold711/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_51_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold70/X fanout327/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X
+ hold400/A fanout57/X m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2
+ fanout240/X hold334/A m_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__a31o_2_B1 m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__and2_2_A/B
+ m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__a2bb2o_2_A1_N/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_buffer\[2\].m_c_buf m_blake2.m_hash256.g_buffer\[2\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[2\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_751 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold770/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR fanout151/A sky130_fd_sc_hd__and4_1
XFILLER_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y
+ fanout224/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_31_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1070 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ hold747/A fanout125/X m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a211o_1
Xhold107 hold107/A VGND VGND VPWR VPWR hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout290/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold129 hold129/A VGND VGND VPWR VPWR hold129/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 hold118/A VGND VGND VPWR VPWR hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout224/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout468/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A/B m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ sky130_fd_sc_hd__xor2_2
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1172/A fanout124/X fanout88/X m_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold840/X fanout543/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout609 fanout610/X VGND VGND VPWR VPWR fanout609/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1030 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold101/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout174/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1170/A hold1103/X fanout586/X VGND VGND VPWR VPWR hold1104/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_S fanout410/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold91/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.res_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_A
+ fanout478/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold158/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout158_A fanout160/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold108/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1097/A
+ fanout604/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__a22o_2_A1 hold769/A fanout291/X
+ fanout279/X hold663/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_40_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__nand2b_2_A_N_A_N
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__mux2_1_A0 hold395/A m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout396/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xhold630 hold630/A VGND VGND VPWR VPWR hold630/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[11\]\[29\]_sky130_fd_sc_hd__o22a_2_A1 hold640/A m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ fanout172/X fanout253/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__o22a_1
Xhold652 hold652/A VGND VGND VPWR VPWR hold652/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold641 hold641/A VGND VGND VPWR VPWR hold641/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 hold663/A VGND VGND VPWR VPWR hold663/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold685 hold685/A VGND VGND VPWR VPWR hold685/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 hold696/A VGND VGND VPWR VPWR hold696/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold674 hold674/A VGND VGND VPWR VPWR hold674/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_49_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_38_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_1
+ fanout418/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR fanout204/A sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A0 hold29/A m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold996/X m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_507 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__a22o_2_A1 hold343/A fanout187/X
+ fanout195/X hold862/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold897/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout26_X fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold748/X fanout562/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_41_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[18\].m_c_buf m_blake2.m_hash256.g_buffer\[18\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[18\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout478/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__a221o_2_B2 hold686/A fanout348/X fanout304/X
+ hold573/A fanout268/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__a221o_2_B2/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_matrix\[3\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__a22o_2_A1 hold604/A fanout190/X
+ fanout198/X hold888/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout291/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ hold542/X VGND VGND VPWR VPWR hold541/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/B
+ sky130_fd_sc_hd__nand3_2
Xm_blake2.m_hash256.m_matrix\[1\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1202/X hold1101/X fanout546/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X data\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1/A2
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_19_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold1043/X m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1031/A sky130_fd_sc_hd__dfxtp_1
Xdata\[3\]_sky130_fd_sc_hd__mux2_1_A1 data\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold7/X
+ fanout600/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_80_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_50_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold760/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout302/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or3_2_A fanout450/X fanout457/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_30_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_65_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold825/X fanout220/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold577/X fanout597/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1 hold987/A fanout348/X
+ fanout260/X m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__and2_2_B fanout428/X hold115/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xfanout439 fanout441/X VGND VGND VPWR VPWR fanout439/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xfanout417 fanout418/X VGND VGND VPWR VPWR fanout417/X sky130_fd_sc_hd__buf_4
Xfanout428 fanout429/X VGND VGND VPWR VPWR fanout428/X sky130_fd_sc_hd__clkbuf_4
Xfanout406 fanout406/A VGND VGND VPWR VPWR fanout406/X sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_18_Left_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_A_N_A_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
XFILLER_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[3\].m_y_buf m_blake2.m_hash256.g_buffer\[3\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[3\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_33_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout275_A fanout276/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[13\]\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold547/X fanout207/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_46_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2
+ fanout274/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout442_A fanout443/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_18_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__or2_2_A hold614/A fanout243/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold954/A fanout59/X fanout71/X hold520/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xfanout35 fanout35/A VGND VGND VPWR VPWR fanout35/X sky130_fd_sc_hd__buf_2
Xfanout46 fanout47/A VGND VGND VPWR VPWR fanout46/X sky130_fd_sc_hd__clkbuf_4
Xfanout24 fanout27/X VGND VGND VPWR VPWR fanout24/X sky130_fd_sc_hd__buf_4
XFILLER_23_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y
+ hold989/A fanout148/X m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y/B1
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/A2
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_11_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout328_X fanout328/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout79 fanout79/A VGND VGND VPWR VPWR fanout79/X sky130_fd_sc_hd__clkbuf_2
Xfanout68 fanout71/A VGND VGND VPWR VPWR fanout68/X sky130_fd_sc_hd__clkbuf_4
Xfanout57 fanout59/A VGND VGND VPWR VPWR fanout57/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold685/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold1204/A fanout132/X fanout141/X hold1041/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__and3_2_A hold244/A fanout465/A fanout373/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold711/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[20\]_sky130_fd_sc_hd__and2_2_X_A fanout354/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold471 hold471/A VGND VGND VPWR VPWR hold471/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__xnor2_2_A hold1054/X m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/X
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xnor2_1
XFILLER_46_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold460 hold460/A VGND VGND VPWR VPWR hold460/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_S fanout213/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold482 hold482/A VGND VGND VPWR VPWR hold482/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold493 hold493/A VGND VGND VPWR VPWR hold493/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1160 hold1160/A VGND VGND VPWR VPWR hold1160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1193 hold1193/A VGND VGND VPWR VPWR hold1193/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1171 hold1171/A VGND VGND VPWR VPWR hold1171/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1182 hold1182/A VGND VGND VPWR VPWR hold1182/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XFILLER_60_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XFILLER_57_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold504/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__a32o_2_A1 hold905/A fanout354/X
+ fanout251/X fanout170/X m_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__a32o_2_A1/X
+ sky130_fd_sc_hd__a32o_1
Xm_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__or2_2_B fanout495/X hold231/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold580/X m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A0 hold24/A m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1088/A fanout26/X fanout50/X m_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout359/X m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ fanout180/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a211o_1
Xclkload16 clkload16/A VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__inv_6
Xm_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR ANTENNA_12/DIODE
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout192/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload27 clkload27/A VGND VGND VPWR VPWR clkload27/Y sky130_fd_sc_hd__inv_12
XTAP_TAPCELL_ROW_11_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold874/X m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout299/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_29_1434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold406/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.fsm_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and4_2_X
+ fanout610/X fanout463/X hold1268/X hash_v_sky130_fd_sc_hd__a211o_2_X/A2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.fsm_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and4_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout31/X fanout39/X
+ hold1177/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_62_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_673 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__or2_2_A hold1239/A fanout391/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_3_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold1215/A fanout35/X m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold958/X hold798/X fanout583/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[19\].m_y_buf m_blake2.m_hash256.g_buffer\[19\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[19\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout233/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_75_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout123/A sky130_fd_sc_hd__and4_1
XFILLER_51_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[15\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold648/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold482/X m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout154/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold413/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold355/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_S fanout203/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout214 fanout216/X VGND VGND VPWR VPWR fanout214/X sky130_fd_sc_hd__buf_6
Xfanout203 fanout204/X VGND VGND VPWR VPWR fanout203/X sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout247 fanout248/X VGND VGND VPWR VPWR fanout247/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout392_A fanout398/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout225 fanout228/A VGND VGND VPWR VPWR fanout225/X sky130_fd_sc_hd__buf_4
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout236 fanout236/A VGND VGND VPWR VPWR fanout236/X sky130_fd_sc_hd__buf_4
Xfanout258 fanout258/A VGND VGND VPWR VPWR fanout258/X sky130_fd_sc_hd__buf_4
XFILLER_59_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout269 fanout269/A VGND VGND VPWR VPWR fanout269/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_31_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_X fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold839/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout278_X fanout278/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[26\]_sky130_fd_sc_hd__o21a_2_A1 hold1267/A fanout367/X
+ fanout169/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[26\]_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold562/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_1
+ fanout413/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR fanout216/A sky130_fd_sc_hd__o21ai_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_data\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold493/X hold1011/A fanout548/X VGND VGND VPWR VPWR hold494/A sky130_fd_sc_hd__mux2_1
XFILLER_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A0 hold72/A m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout518/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__a311o_2_A1_A2 fanout354/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold705/X hold641/X fanout605/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B1
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__or2_2_B fanout498/X hold18/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[6\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1093/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_46_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold290 hold290/A VGND VGND VPWR VPWR hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1146/X m_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout541/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_827 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout17/X hold675/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[22\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/X m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1 fanout461/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/C m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/X
+ sky130_fd_sc_hd__o31a_1
Xm_blake2.m_hash256.m_matrix\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1151/X m_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout581/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_53_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/B2 hold1041/X fanout569/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_C_sky130_fd_sc_hd__o31a_2_X_A1
+ fanout407/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1/Y m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1/X
+ VGND VGND VPWR VPWR fanout224/A sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold746/X fanout329/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_702 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_B m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2
+ fanout285/X m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2/X
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_S fanout224/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B fanout487/X hold121/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_A1 m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_2
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XFILLER_9_1336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[10\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold541/X hold1236/A fanout566/X VGND VGND VPWR VPWR hold542/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/A
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/B
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ sky130_fd_sc_hd__and3_1
Xinput3 ui_in[0] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[30\].m_y_buf m_blake2.m_hash256.g_buffer\[30\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[30\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B fanout484/X hold140/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout238_A fanout239/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold218/X fanout166/X m_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout405_A fanout406/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/D
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A1 VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[29\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout170/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout403/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__o21ai_2_A1 hold578/A fanout368/X
+ fanout193/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__a21oi_2_A1_A2 fanout282/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__xnor2_2_A hold401/A hold822/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XFILLER_47_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout87/A sky130_fd_sc_hd__and4_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_io.m_config.ll_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X hold1258/X
+ VGND VGND VPWR VPWR hold255/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X_A1 fanout182/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold203/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_687 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold443/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__or2_2_A hold642/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold1022/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B fanout484/X hold80/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_io.m_block_data.data_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ ena_sky130_fd_sc_hd__or2_2_B/A m_io.m_block_data.data_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold1263/X fanout335/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhash\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hash\[7\]_sky130_fd_sc_hd__and2_2_B/B fanout335/X VGND VGND VPWR VPWR hash\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout343/X m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__a22o_2_A1 hold465/A fanout291/X
+ fanout406/X hold770/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR fanout75/A sky130_fd_sc_hd__nor2_2
XFILLER_26_1415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__a31o_2_B1 ANTENNA_11/DIODE
+ m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__and2_2_A/B
+ m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X m_blake2.m_hash256.g_buffer\[2\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout193/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.fsm_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C
+ m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout155/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_S fanout300/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__mux2_1_A0 hold1221/A m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout532/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_io.m_config.ll_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold196/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1
+ fanout197/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout527/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2/X
+ m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout403/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout193/X m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout176/X fanout270/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__xnor2_2_A hold450/A hold759/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2 m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ fanout259/X fanout304/X m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__or2_2_A/A m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/C1
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/X sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N_X m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N/Y
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N/X
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1/X
+ sky130_fd_sc_hd__o21ba_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1197/X hold1158/X fanout604/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout188_A fanout189/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C fanout249/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout176/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout355_A fanout361/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold183/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_4
XTAP_TAPCELL_ROW_23_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout522_A fanout524/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ hold352/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold1012/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout408_X fanout408/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1 hold1218/A fanout343/X
+ fanout259/X m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold754/X m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout418/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_S fanout213/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__xnor2_2_A hold245/A hold738/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1206/X
+ fanout562/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_7_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_2
XFILLER_56_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout56_X fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_963 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A0 hold84/A m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ hold1240/A fanout307/X m_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
XFILLER_44_911 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_6_Left_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout413/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold844/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1
+ fanout287/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__xnor2_2_A hold828/A hold823/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout66/X
+ fanout79/X hold983/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout170/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A0 hold219/A m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/C sky130_fd_sc_hd__and2_1
XFILLER_8_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1162/X m_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout549/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__or2_2_B fanout488/X hold167/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[14\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold717/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout288/X m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout295/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1033/A fanout50/X fanout46/X hold1096/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout416/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold249/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__xnor2_2_A hold1212/A hold1048/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_54_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold1186/A fanout91/X m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout107/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_35_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold606/X fanout588/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[5\]_sky130_fd_sc_hd__mux2_1_A1_A1 hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhold801 hold801/A VGND VGND VPWR VPWR hold801/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold812 hold812/A VGND VGND VPWR VPWR hold812/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 hold823/A VGND VGND VPWR VPWR hold823/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold845 hold845/A VGND VGND VPWR VPWR hold845/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold834 hold834/A VGND VGND VPWR VPWR hold834/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_S fanout204/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xhold878 hold878/A VGND VGND VPWR VPWR hold878/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold856 hold856/A VGND VGND VPWR VPWR hold856/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 hold889/A VGND VGND VPWR VPWR hold889/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 hold867/A VGND VGND VPWR VPWR hold867/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout425/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout26/X fanout78/X
+ m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_51_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout472_A fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout417/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A0 hold222/A m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout511/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout260_X fanout260/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__xnor2_2_A hold302/A hold1219/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold185/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1161/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/X m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X/A1
+ sky130_fd_sc_hd__nand2b_1
Xm_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A/B sky130_fd_sc_hd__xor2_4
XFILLER_26_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ hold1141/X VGND VGND VPWR VPWR hold1140/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__or2_2_B fanout487/X hold62/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X
+ m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_21_693 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2_C_sky130_fd_sc_hd__or2_2_X
+ fanout457/X fanout459/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/C
+ sky130_fd_sc_hd__or2_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout193/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold698/A fanout58/X fanout47/X hold571/A m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__and2b_2_B m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1/B1 sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout404/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ hold750/A fanout33/X m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a211o_1
XFILLER_76_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21boi_2_Y
+ hold652/A m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__o311a_2_A1/X VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21boi_1
Xm_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0_A1_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C/X
+ m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0_A1_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold750/A fanout125/X fanout85/X m_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_1180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_B
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout89/X
+ fanout145/X hold896/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_A
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.g_buffer\[6\].m_c_buf m_blake2.m_hash256.g_buffer\[6\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[6\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2
+ fanout487/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A/Y fanout274/X
+ m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/X
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B fanout490/X hold110/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__a22o_2_A1 hold689/A m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__or3_2_B/X fanout249/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/B2 sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold108 hold108/A VGND VGND VPWR VPWR hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold924/X hold1193/A fanout596/X VGND VGND VPWR VPWR hold925/A sky130_fd_sc_hd__mux2_1
Xhold119 hold119/A VGND VGND VPWR VPWR hold119/X sky130_fd_sc_hd__dlygate4sd3_1
Xena_sky130_fd_sc_hd__or2_2_B ena_sky130_fd_sc_hd__or2_2_B/A input1/X VGND VGND VPWR
+ VPWR ena_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_S fanout224/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_io.en_q_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A ena_sky130_fd_sc_hd__or2_2_B/X VGND
+ VGND VPWR VPWR fanout1/A sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold696/A fanout34/X fanout46/X hold1133/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_39_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X
+ fanout191/X m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__nand2_2_B/Y
+ fanout274/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_50_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold352/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold902/A fanout26/X fanout82/X hold1031/A m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_40_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout318_A fanout323/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout220_A fanout220/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold620 hold620/A VGND VGND VPWR VPWR hold620/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
Xhold642 hold642/A VGND VGND VPWR VPWR hold642/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout106_X fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold631 hold631/A VGND VGND VPWR VPWR hold631/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold653 hold653/A VGND VGND VPWR VPWR hold653/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold686 hold686/A VGND VGND VPWR VPWR hold686/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 hold664/A VGND VGND VPWR VPWR hold664/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 hold697/A VGND VGND VPWR VPWR hold697/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold675 hold675/A VGND VGND VPWR VPWR hold675/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X
+ data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/X m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ fanout611/X m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A hold523/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_38_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold230/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold989/X hold1156/A fanout548/X VGND VGND VPWR VPWR hold990/A sky130_fd_sc_hd__mux2_1
XFILLER_57_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1128/X fanout226/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold29/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__nand2_2_B fanout440/X hold181/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold193/X fanout605/X
+ VGND VGND VPWR VPWR hold194/A sky130_fd_sc_hd__mux2_1
XFILLER_60_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[13\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[13\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold497/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__a21o_2_A1 hold19/X fanout319/X
+ m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__nor2_2_B fanout497/X hold104/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_14_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ hold1260/X m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout426/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.m_matrix\[13\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[13\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1029/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_20_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_20_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_2
Xm_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold153/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[12\]\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1083/X fanout226/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold375/A m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout363/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A2/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o21a_2_A2/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B/X
+ sky130_fd_sc_hd__or4_1
Xm_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a31o_2_X
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A3 m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B
+ m_io.cmd\[2\]_sky130_fd_sc_hd__nor2_2_A/Y m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/A
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_68_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1_sky130_fd_sc_hd__a21o_2_A2
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/B1
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1_sky130_fd_sc_hd__a21o_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B/A
+ sky130_fd_sc_hd__a21o_1
XFILLER_27_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold48/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_75_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A0 hold40/A m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold226/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold241/X m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout236/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout406/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold637/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold282/X m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_9_Left_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/X sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_80_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_11_clk clkload1/A VGND VGND VPWR VPWR clkload17/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1 m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__a22o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__xor2_2_A hold292/A hold473/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__a31o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1/X m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_30_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/B2
+ hold486/X fanout557/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__a22o_2_A1 hold471/A fanout192/X
+ fanout200/X hold855/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[10\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold962/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold1017/X m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout177/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout407 fanout408/A VGND VGND VPWR VPWR fanout407/X sky130_fd_sc_hd__buf_6
Xfanout418 fanout420/A VGND VGND VPWR VPWR fanout418/X sky130_fd_sc_hd__buf_4
Xfanout429 fanout431/X VGND VGND VPWR VPWR fanout429/X sky130_fd_sc_hd__buf_2
XFILLER_80_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_blake2.m_hash256.g_buffer\[2\].m_y_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_buffer\[7\].m_y_buf m_blake2.m_hash256.g_buffer\[7\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[7\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout268_A fanout269/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout287/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_A
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout210/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1176/A sky130_fd_sc_hd__dfxtp_1
Xfanout47 fanout47/A VGND VGND VPWR VPWR fanout47/X sky130_fd_sc_hd__clkbuf_2
XFILLER_35_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout25 fanout27/X VGND VGND VPWR VPWR fanout25/X sky130_fd_sc_hd__buf_2
XFILLER_23_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout36 fanout39/A VGND VGND VPWR VPWR fanout36/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout435_A fanout443/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold402/A m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout397/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xfanout58 fanout59/A VGND VGND VPWR VPWR fanout58/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xfanout69 fanout71/A VGND VGND VPWR VPWR fanout69/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_939 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B fanout488/X hold34/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_52_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout223_X fanout223/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X fanout1/X
+ fanout609/X input11/X VGND VGND VPWR VPWR m_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold461 hold461/A VGND VGND VPWR VPWR hold461/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 hold472/A VGND VGND VPWR VPWR hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 hold450/A VGND VGND VPWR VPWR hold450/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 hold483/A VGND VGND VPWR VPWR hold483/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[13\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1011/X hold959/X fanout548/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold494 hold494/A VGND VGND VPWR VPWR hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A fanout83/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_69_clk clkload0/A VGND VGND VPWR VPWR clkbuf_leaf_69_clk/X sky130_fd_sc_hd__clkbuf_8
Xhold1150 hold1150/A VGND VGND VPWR VPWR hold1150/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_674 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold978/X fanout206/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/C fanout424/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
Xhold1161 hold1161/A VGND VGND VPWR VPWR hold1161/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[14\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1072/X m_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout595/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold1194 hold1194/A VGND VGND VPWR VPWR hold1194/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[10\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold764/X hold994/A fanout585/X VGND VGND VPWR VPWR hold765/A sky130_fd_sc_hd__mux2_1
Xhold1183 hold1183/A VGND VGND VPWR VPWR hold1183/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[1\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[1\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold772/A sky130_fd_sc_hd__dfxtp_1
Xhold1172 hold1172/A VGND VGND VPWR VPWR hold1172/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
XFILLER_73_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold62/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_880 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A1 m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_0_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout256/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1198/A fanout58/X fanout46/X hold1095/A m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold24/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold800/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout349/X m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X fanout256/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload17 clkload17/A VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__inv_8
Xm_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold234/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X m_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold77/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_983 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload28 clkload28/A VGND VGND VPWR VPWR clkload28/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold870/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[3\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold937/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__o22a_2_A2/X
+ hold143/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold593/X fanout204/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/A
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/X m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2/A2_N
+ m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout178/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout183/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_0_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_0_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__a31o_2_B1_A3
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold776/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[11\]\[31\]_sky130_fd_sc_hd__or2_2_A hold1182/A fanout388/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[31\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__a211oi_2_A1 hold779/A fanout402/X
+ m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__a22o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__a211oi_2_A1/Y
+ sky130_fd_sc_hd__a211oi_1
Xm_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold859/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[5\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[5\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold328/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.g_buffer\[10\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_17_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A hold315/A hold844/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A0 hold175/A m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout508/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout621/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__mux2_1_A0 hold109/A m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A_B fanout485/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold328/A fanout112/X m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XFILLER_69_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout260/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold319/X hold445/X fanout606/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1140/X fanout591/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout204 fanout204/A VGND VGND VPWR VPWR fanout204/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[7\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold780/A sky130_fd_sc_hd__dfxtp_1
Xfanout226 fanout228/A VGND VGND VPWR VPWR fanout226/X sky130_fd_sc_hd__buf_2
Xfanout237 fanout239/A VGND VGND VPWR VPWR fanout237/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_matrix\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold782/X VGND VGND VPWR VPWR hold781/A sky130_fd_sc_hd__dfxtp_1
Xfanout215 fanout216/X VGND VGND VPWR VPWR fanout215/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xfanout248 fanout248/A VGND VGND VPWR VPWR fanout248/X sky130_fd_sc_hd__clkbuf_2
Xfanout259 fanout260/X VGND VGND VPWR VPWR fanout259/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout385_A fanout399/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X hold185/A m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/A2
+ m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/B1 VGND VGND VPWR VPWR uio_out_sky130_fd_sc_hd__buf_2_X/A
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__a21o_2_B1 m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/C m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_54_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__a21o_2_X/A2
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/C sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout173_X fanout173/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout278/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_59_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_65_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[9\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold680/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold72/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__a311o_2_A1_A3 fanout249/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold421/X fanout563/X
+ VGND VGND VPWR VPWR hold422/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__xor2_2_A hold627/A hold189/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold280 hold280/A VGND VGND VPWR VPWR hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold291 hold291/A VGND VGND VPWR VPWR hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout86_X fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout197/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__and2_2_B fanout430/X hold101/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_63_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_config.ll_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X m_io.m_config.ll_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold303/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_64_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout119/A sky130_fd_sc_hd__and4_2
XFILLER_46_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2 fanout458/X fanout461/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2/X
+ sky130_fd_sc_hd__o31a_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__o21a_2_A1_A2 fanout385/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A0 hold187/A m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout529/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_B2
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout420/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/B sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_75_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_17_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold929/X hold911/X fanout597/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B/A
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_B2_sky130_fd_sc_hd__inv_2_Y
+ hold1162/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/B2
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout200/X m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout192/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xinput4 ui_in[1] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_65_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__and2_2_B_A fanout434/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A/C
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2_X m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y
+ m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__o21ai_2
XFILLER_25_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B
+ fanout266/X m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_75_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[9\]_sky130_fd_sc_hd__or2_2_A hold528/A fanout241/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[9\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/B1
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/A3
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_A
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21oi_2_B1_A1
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__or2_2_B_A fanout500/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout300_A fanout301/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold735/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_905 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_A
+ fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XFILLER_0_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout290_X fanout290/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout394/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_56_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or3b_2_B/X
+ m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
XFILLER_27_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_67_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand2_2_B
+ fanout471/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR fanout274/A sky130_fd_sc_hd__nand2_8
XANTENNA_fanout46_A fanout47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A0 hold111/A m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout518/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold662/A fanout109/X fanout145/X m_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1
+ fanout407/X m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND
+ VGND VPWR VPWR fanout252/A sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_26_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold123/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_io.m_block_data.data_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_block_data.data_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/B
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_io.m_block_data.data_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and3b_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/A
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/Y
+ sky130_fd_sc_hd__nand3_2
Xm_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0 m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y
+ hold77/A fanout430/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0 hold583/X m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout534/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B_B m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout590 fanout608/X VGND VGND VPWR VPWR fanout590/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_matrix\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1151/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_931 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_B1
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xblock_first_sky130_fd_sc_hd__a32o_2_B2 block_first_sky130_fd_sc_hd__a32o_2_B2/A1
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A2 block_last_sky130_fd_sc_hd__a32o_2_B2/A3
+ block_last_sky130_fd_sc_hd__a32o_2_B2/B1 hold13/A VGND VGND VPWR VPWR block_first_sky130_fd_sc_hd__a32o_2_B2/X
+ sky130_fd_sc_hd__a32o_1
Xm_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[2\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold936/X hold881/X fanout598/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold1216/X fanout221/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_72_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__a22o_2_A1 hold23/X fanout338/X
+ m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_77_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__or2_2_A hold573/A fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X hold583/X fanout275/X m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/C1 m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/D1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/X sky130_fd_sc_hd__a2111o_1
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_A2_sky130_fd_sc_hd__and2_2_X
+ fanout355/X fanout253/X VGND VGND VPWR VPWR fanout174/A sky130_fd_sc_hd__and2_2
Xm_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X
+ fanout269/A m_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__and4_1
Xm_blake2.m_hash256.m_matrix\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold739/X hold646/X fanout588/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[13\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout181/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2_X_sky130_fd_sc_hd__o21a_2_A2
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/C m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/C
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1 hold514/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout425/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.m_matrix\[9\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1172/X hold1188/A fanout541/X VGND VGND VPWR VPWR hold1173/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__a31o_2_B1 m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__and2_2_A/B
+ m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
Xm_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1109/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__mux2_1_A1_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_975 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold415/X hold328/X fanout542/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_52_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__xnor2_2_B hold1267/A hold510/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout250_A fanout252/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout348_A fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ sky130_fd_sc_hd__nor2_1
XFILLER_80_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout269/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1133/X hold1095/X fanout554/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_2
XANTENNA_fanout136_X fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__xnor2_2_A hold355/A hold1091/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1040/X
+ fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout303_X fanout303/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_matrix\[0\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold453/X m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout605/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__mux2_1_A0_A0 m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold63/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_S fanout412/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_768 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_7_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/X fanout609/X input9/X VGND VGND VPWR VPWR m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
XFILLER_48_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_29_975 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold84/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__and3_2_C fanout448/X fanout479/X
+ hold95/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XFILLER_44_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold861/A fanout30/X fanout54/X m_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A_1 fanout472/X fanout407/X
+ VGND VGND VPWR VPWR fanout295/A sky130_fd_sc_hd__nor2_2
XFILLER_19_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1008 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold219/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y hash\[0\]_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0_A1_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__nor2_2_B fanout483/X hold180/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_7_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__nor2_2_B_A fanout497/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_B1
+ fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold244/X fanout162/X m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold779/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_c_buf\[0\]_sky130_fd_sc_hd__a211o_2_X m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.g_c_buf\[0\]_sky130_fd_sc_hd__a211o_2_X/A2 m_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__o21a_2_A1/X
+ m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__o21a_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[0\].m_c_buf/A sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold257/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout171/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout252/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__mux2_1_A0 hold105/A m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_17_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N_A1
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_33_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold589/A fanout127/X m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout107/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout90/X fanout138/X
+ hold1095/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[28\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold802 hold802/A VGND VGND VPWR VPWR hold802/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__xnor2_2_B hold991/A hold751/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold824 hold824/A VGND VGND VPWR VPWR hold824/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold813 hold813/A VGND VGND VPWR VPWR hold813/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 hold846/A VGND VGND VPWR VPWR hold846/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold835 hold835/A VGND VGND VPWR VPWR hold835/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold857 hold857/A VGND VGND VPWR VPWR hold857/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold868 hold868/A VGND VGND VPWR VPWR hold868/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 hold879/A VGND VGND VPWR VPWR hold879/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_44_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout298_A fanout299/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold74/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_S fanout371/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout465_A fanout465/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_28_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold222/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D_sky130_fd_sc_hd__a22o_2_X_B2 hash\[6\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D_sky130_fd_sc_hd__a22o_2_X_A1 m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold725/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__a22o_2_A1 hold287/A fanout289/X
+ fanout284/X hold327/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_77_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__inv_2_Y
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X/B1
+ sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_49_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout420_X fanout420/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__o22a_2_A1_B1 fanout173/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A/B
+ fanout358/X fanout262/X hold1255/A m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[13\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold861/X m_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout595/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A0 hold170/A m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout536/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
XFILLER_62_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__a22o_2_A1 hold673/A fanout191/X
+ fanout199/X hold661/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__a32o_2_A1 m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/A
+ fanout345/X fanout250/X fanout171/X m_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__a32o_2_A1/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_5_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_731 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_934 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout182/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1254/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__a22o_2_A1 hold517/A fanout188/X
+ fanout196/X hold804/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_32_959 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ hold255/X fanout304/X m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y/B sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_S fanout208/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold350/X m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_C_sky130_fd_sc_hd__o31a_2_X
+ fanout458/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/D
+ fanout444/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_8_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold109 hold109/A VGND VGND VPWR VPWR hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_S fanout215/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X data\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold239/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold344/X m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout301/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1_sky130_fd_sc_hd__or2_2_X
+ hold483/A fanout102/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A1
+ sky130_fd_sc_hd__or2_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1 hold1241/A fanout343/X
+ fanout259/X m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold916/A sky130_fd_sc_hd__dfxtp_1
Xm_io.cmd\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X m_io.cmd\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__a32o_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_54_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold649/X m_blake2.m_hash256.m_matrix\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout606/X
+ VGND VGND VPWR VPWR hold650/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1265/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_22_Left_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_40_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout213_A fanout216/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold610 hold610/A VGND VGND VPWR VPWR hold610/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout195/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold737/A sky130_fd_sc_hd__dfxtp_1
Xhold621 hold621/A VGND VGND VPWR VPWR hold621/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold643 hold643/A VGND VGND VPWR VPWR hold643/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 hold632/A VGND VGND VPWR VPWR hold632/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_31_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold654 hold654/A VGND VGND VPWR VPWR hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_9_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold687 hold687/A VGND VGND VPWR VPWR hold687/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 hold676/A VGND VGND VPWR VPWR hold676/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 hold665/A VGND VGND VPWR VPWR hold665/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold987/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold698 hold698/A VGND VGND VPWR VPWR hold698/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold489/X m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/A fanout263/X
+ m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__a221o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_1
XFILLER_58_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2
+ fanout292/X m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2/X
+ sky130_fd_sc_hd__a21bo_1
Xm_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold806/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X/A
+ sky130_fd_sc_hd__xnor2_1
XFILLER_41_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A hold579/A fanout354/X
+ fanout249/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XFILLER_16_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_c_buf\[8\]_sky130_fd_sc_hd__a211o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold681/X m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1021 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold375/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold493/A fanout80/X m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[10\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold470/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold478/X m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout184/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold558/A fanout129/X fanout117/X hold1199/A m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout229/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold40/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold734/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_19_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__nand2_2_B fanout439/X hold124/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__a211oi_2_A1 hold460/A fanout280/X
+ m_blake2.m_hash256.v_q\[1\]\[27\]_sky130_fd_sc_hd__a22o_2_A1/X fanout390/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__a211oi_2_A1/Y
+ sky130_fd_sc_hd__a211oi_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout90/X
+ fanout146/X hold912/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_80_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold595/X m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold749/X hold638/X fanout589/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1117/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ hold236/X VGND VGND VPWR VPWR hold235/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__a22o_2_A1_B2 fanout252/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2 fanout451/X fanout454/X
+ fanout460/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/D m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/X
+ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_30_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout594/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold271/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1145/X fanout227/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.g_c_buf\[27\]_sky130_fd_sc_hd__o22a_2_X hold1191/A fanout175/A
+ m_blake2.m_hash256.g_c_buf\[27\]_sky130_fd_sc_hd__o22a_2_X/B1 m_blake2.m_hash256.g_c_buf\[27\]_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[27\].m_c_buf/A sky130_fd_sc_hd__o22a_1
XFILLER_28_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout419 fanout420/X VGND VGND VPWR VPWR fanout419/X sky130_fd_sc_hd__buf_4
XFILLER_28_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout408 fanout408/A VGND VGND VPWR VPWR fanout408/X sky130_fd_sc_hd__buf_2
XFILLER_80_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_2
Xm_blake2.m_hash256.m_matrix\[15\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ data\[2\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_804 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[14\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold387/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout405/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A2
+ sky130_fd_sc_hd__a22o_2
XFILLER_55_837 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold1044/X m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout153/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout163_A fanout168/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold404/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout26 fanout27/X VGND VGND VPWR VPWR fanout26/X sky130_fd_sc_hd__clkbuf_4
XFILLER_39_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout110/X
+ fanout142/X hold1192/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xfanout37 fanout39/A VGND VGND VPWR VPWR fanout37/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout330_A fanout342/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout59 fanout59/A VGND VGND VPWR VPWR fanout59/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2/X
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout428_A fanout429/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout48 fanout51/A VGND VGND VPWR VPWR fanout48/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold402/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/A
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout216_X fanout216/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[14\]_sky130_fd_sc_hd__mux2_1_A1_S fanout223/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold451 hold451/A VGND VGND VPWR VPWR hold451/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold440 hold440/A VGND VGND VPWR VPWR hold440/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 hold462/A VGND VGND VPWR VPWR hold462/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 hold495/A VGND VGND VPWR VPWR hold495/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 hold484/A VGND VGND VPWR VPWR hold484/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xhold473 hold473/A VGND VGND VPWR VPWR hold473/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[8\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold682/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1 fanout449/X fanout450/X
+ fanout453/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hash\[0\]_sky130_fd_sc_hd__or2_2_B_B hash\[0\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1140 hold1140/A VGND VGND VPWR VPWR hold1140/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/C
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/X
+ sky130_fd_sc_hd__or4_1
Xhold1151 hold1151/A VGND VGND VPWR VPWR hold1151/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_2
Xm_blake2.m_hash256.v_q\[8\]\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1035/X fanout223/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1184 hold1184/A VGND VGND VPWR VPWR hold1184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1173 hold1173/A VGND VGND VPWR VPWR hold1173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1162 hold1162/A VGND VGND VPWR VPWR hold1162/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
Xhold1195 hold1195/A VGND VGND VPWR VPWR hold1195/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2
+ m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__a211oi_2_A1/Y m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2/Y
+ fanout405/X m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ sky130_fd_sc_hd__a2bb2o_2
XTAP_TAPCELL_ROW_0_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.m_matrix\[6\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1209/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
Xclkload18 clkload18/A VGND VGND VPWR VPWR clkload18/X sky130_fd_sc_hd__clkbuf_8
Xclkload29 clkload29/A VGND VGND VPWR VPWR clkload29/Y sky130_fd_sc_hd__clkinv_2
XFILLER_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_11_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A1_N
+ fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1088/X m_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout591/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[8\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ hold647/X VGND VGND VPWR VPWR hold646/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_63_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B/B sky130_fd_sc_hd__dfxtp_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__or2_2_B_A fanout485/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_60_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold175/X fanout317/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold109/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold856/A hold407/X fanout540/X VGND VGND VPWR VPWR hold408/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1/A1
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__o31a_2_A2 fanout408/X m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/A
+ fanout388/X fanout249/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[27\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__o31a_1
Xfanout205 fanout208/X VGND VGND VPWR VPWR fanout205/X sky130_fd_sc_hd__buf_4
Xm_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout241/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout216 fanout216/A VGND VGND VPWR VPWR fanout216/X sky130_fd_sc_hd__buf_4
Xfanout227 fanout228/X VGND VGND VPWR VPWR fanout227/X sky130_fd_sc_hd__buf_4
Xfanout238 fanout239/X VGND VGND VPWR VPWR fanout238/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_B1
+ fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout249 fanout249/A VGND VGND VPWR VPWR fanout249/X sky130_fd_sc_hd__buf_6
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/A1
+ sky130_fd_sc_hd__nand2_1
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout280_A fanout282/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ sky130_fd_sc_hd__and2b_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout300/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_884 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_704 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A0 hold153/A m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1074/A fanout42/X fanout78/X m_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_B2
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout500_X fanout500/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__xnor2_2_A hold395/A hold1092/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A0 hold104/A m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold270 hold270/A VGND VGND VPWR VPWR hold270/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ hold1028/X VGND VGND VPWR VPWR hold1027/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout426/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
Xhold281 hold281/A VGND VGND VPWR VPWR hold281/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold292 hold292/A VGND VGND VPWR VPWR hold292/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__or2_1
XFILLER_77_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X hold351/A fanout18/X m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[25\].m_y_buf/A sky130_fd_sc_hd__o22a_1
XFILLER_74_910 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B/B sky130_fd_sc_hd__dfxtp_1
XFILLER_24_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout30/X fanout74/X
+ hold988/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_46_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout115/A sky130_fd_sc_hd__and4_2
Xm_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold178/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A1_S fanout341/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout100/X m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o32a_4
Xm_blake2.m_hash256.m_matrix\[9\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1188/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_Y
+ fanout400/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__a22o_2_A1 hold438/A fanout289/X
+ fanout277/X hold481/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold187/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_A
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout583/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A0_S fanout520/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_75_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_S fanout213/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_71_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_71_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.g_buffer\[7\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/B m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2
+ fanout240/A hold986/A m_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XFILLER_9_1316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1 m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_matrix\[11\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1040/X m_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout542/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__and2_2_B fanout439/X hold58/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xinput5 ui_in[2] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.g_idx_next\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ fanout474/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B
+ sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold797/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout66/X fanout42/X
+ m_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout413/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_998 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_80_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout446/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/A1
+ sky130_fd_sc_hd__inv_2
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ sky130_fd_sc_hd__a21bo_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold232/A m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__or2_2_B/X fanout392/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_33_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold72/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_20_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_60_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y
+ fanout51/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout126_A fanout127/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1038/A fanout57/X fanout25/X hold897/A m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ hold1199/A fanout29/X m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21bo_2_X
+ m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout495_A fanout497/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout283_X fanout283/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold148/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold743/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1017 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_67_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C/A
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/A1
+ sky130_fd_sc_hd__a21oi_4
Xm_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold111/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_35_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout275/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout595/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout39_A fanout39/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_26_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_S fanout203/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold660/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold601/X hold944/A fanout592/X VGND VGND VPWR VPWR hold602/A sky130_fd_sc_hd__mux2_1
XFILLER_65_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.g_buffer\[13\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__and2_2_B fanout431/X hold42/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_66_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout591 fanout592/X VGND VGND VPWR VPWR fanout591/X sky130_fd_sc_hd__clkbuf_4
Xfanout580 fanout582/X VGND VGND VPWR VPWR fanout580/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1_A2 fanout377/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A0 hold205/A m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout528/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout420/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_61_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout80/X
+ fanout64/X hold613/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_467 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2
+ fanout284/X m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout277/X fanout346/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or4_2_A fanout454/X fanout457/X
+ fanout459/X fanout461/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_A
+ fanout413/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_78_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_77_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__xnor2_2_A hold326/A hold1128/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[10\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold656/X hold1076/A fanout606/X VGND VGND VPWR VPWR hold657/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XFILLER_29_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2_A1 m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2
+ fanout189/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout196/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y fanout271/X m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ hold1261/X m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ fanout423/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_62_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout243_A fanout248/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__xnor2_2_A hold482/A hold769/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_10 fanout170/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout410_A fanout412/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout508_A fanout509/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_S fanout223/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_63_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B fanout490/X hold144/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_7_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.fsm_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.fsm_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash_v_sky130_fd_sc_hd__a211o_2_X/A2 sky130_fd_sc_hd__dfxtp_1
XFILLER_60_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ ANTENNA_11/DIODE m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XFILLER_46_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout316/X VGND VGND VPWR VPWR hash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A2
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_16_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout157/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__mux2_1_A1_S fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold19/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21boi_2_B1_N
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1/Y m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1/B1
+ sky130_fd_sc_hd__a21boi_1
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold624/X hold668/A fanout601/X VGND VGND VPWR VPWR hold625/A sky130_fd_sc_hd__mux2_1
XFILLER_46_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold594/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout196/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout188/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold294/A m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__and2_2_B/X fanout397/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N_A2
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold397/A fanout27/X fanout31/X hold1099/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold803 hold803/A VGND VGND VPWR VPWR hold803/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 hold836/A VGND VGND VPWR VPWR hold836/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 hold814/A VGND VGND VPWR VPWR hold814/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 hold825/A VGND VGND VPWR VPWR hold825/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold847 hold847/A VGND VGND VPWR VPWR hold847/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold858 hold858/A VGND VGND VPWR VPWR hold858/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 hold869/A VGND VGND VPWR VPWR hold869/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold724/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout198/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout193_A fanout194/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[13\]\[3\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold809/X fanout207/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold579/X m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout155/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout360_A fanout361/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold270/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_787 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__o21a_2_A1 hold1220/A fanout370/X
+ fanout254/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__o22a_2_A1_B2 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout413_X fanout413/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1189/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold331/X fanout603/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1030/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_B1
+ fanout350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold170/X fanout340/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1120/X m_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout580/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[13\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold748/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout404/X m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_2
XFILLER_5_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1050/X hold1026/A fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_1238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__a22o_2_A1 hold480/A fanout292/X
+ fanout286/X hold442/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_21_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_56_1229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A
+ fanout499/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__and2_2_B_A fanout430/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__or2_2_A hold263/A fanout383/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_44_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold26/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XANTENNA_data\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1266/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold405/A m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout389/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2 m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A2 m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ sky130_fd_sc_hd__a22oi_1
Xm_blake2.m_hash256.m_matrix\[0\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/B2 hold1001/X fanout598/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__mux2_1_A0 hold215/A m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout516/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold1267/X m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold1139/X m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout413/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xdata\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold179/X fanout308/X VGND VGND VPWR VPWR data\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1045/X fanout540/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N/X
+ sky130_fd_sc_hd__or3b_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X/A
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__a22o_2_A1 hold297/A fanout187/X
+ fanout195/X hold972/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2 m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ fanout357/X fanout306/X hold461/A fanout269/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2/X
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_44_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[12\]\[18\]_sky130_fd_sc_hd__nand2_2_A hold636/A fanout347/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/C1 sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_44_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold266/X m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1112/A fanout41/X fanout77/X hold564/A m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout206_A fanout207/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold611 hold611/A VGND VGND VPWR VPWR hold611/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold769/A sky130_fd_sc_hd__dfxtp_1
Xhold600 hold600/A VGND VGND VPWR VPWR hold600/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold622 hold622/A VGND VGND VPWR VPWR hold622/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 hold644/A VGND VGND VPWR VPWR hold644/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 hold633/A VGND VGND VPWR VPWR hold633/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A_Y fanout406/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold655 hold655/A VGND VGND VPWR VPWR hold655/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.g_buffer\[7\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xhold666 hold666/A VGND VGND VPWR VPWR hold666/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 hold677/A VGND VGND VPWR VPWR hold677/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 hold688/A VGND VGND VPWR VPWR hold688/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold699 hold699/A VGND VGND VPWR VPWR hold699/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/B m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/B
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold823/X m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout196_X fanout196/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XFILLER_57_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold609/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__and2b_2_B fanout466/X fanout462/X
+ VGND VGND VPWR VPWR fanout399/A sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold658/A fanout118/X fanout98/X m_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[11\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[11\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold304/A m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout373/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold306/X fanout162/X m_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold447/X fanout218/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold688/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_A1
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_B2
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B/B
+ m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout523/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold16/X fanout598/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold343/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2
+ m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/A3
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout196/X m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout188/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[14\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold515/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.v_q\[13\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold285/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__a22o_2_A1_B2 fanout408/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__a211o_2_A1 hold1014/A fanout278/X
+ m_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__a22o_2_A1/X fanout363/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.m_matrix\[1\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ hold903/X VGND VGND VPWR VPWR hold902/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1181/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold604/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold795/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout251/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout291/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_29_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold578/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold872/X fanout220/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_32_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[3\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1057/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold231/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1157/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold449/X m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout418/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout174/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A hold318/A fanout288/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_4
Xm_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold875/X fanout204/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold147/X fanout310/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout162/X m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout616/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_28_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR hold829/A sky130_fd_sc_hd__dfxtp_1
Xfanout409 fanout410/X VGND VGND VPWR VPWR fanout409/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold426/X m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout160/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold749/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold721/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2/Y
+ m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/A2
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.g_buffer\[15\].m_c_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ fanout358/X fanout262/X m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__and3_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_66_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.m_matrix\[11\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1063/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_54_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__and3_2_B_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout57/X fanout36/X
+ hold1070/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A0 hold198/A m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout518/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/B m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout126/X fanout142/X
+ hold1001/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X/D1
+ sky130_fd_sc_hd__a22o_1
Xfanout27 fanout27/A VGND VGND VPWR VPWR fanout27/X sky130_fd_sc_hd__buf_2
Xfanout38 fanout39/A VGND VGND VPWR VPWR fanout38/X sky130_fd_sc_hd__clkbuf_4
Xfanout16 fanout19/A VGND VGND VPWR VPWR fanout16/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout156_A fanout156/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout65/X
+ fanout76/X hold950/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xfanout49 fanout51/A VGND VGND VPWR VPWR fanout49/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_matrix\[13\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[13\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1199/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout323_A fanout342/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__a22o_2_A1_A1 m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ hold521/X VGND VGND VPWR VPWR hold520/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold59/A m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout530/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ hold552/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold570/X m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout239/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_X fanout209/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold452 hold452/A VGND VGND VPWR VPWR hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 hold430/A VGND VGND VPWR VPWR hold430/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 hold441/A VGND VGND VPWR VPWR hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 hold463/A VGND VGND VPWR VPWR hold463/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold474 hold474/A VGND VGND VPWR VPWR hold474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 hold485/A VGND VGND VPWR VPWR hold485/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y
+ fanout473/X fanout477/X VGND VGND VPWR VPWR fanout400/A sky130_fd_sc_hd__nand2_2
Xhold496 hold496/A VGND VGND VPWR VPWR hold496/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout480_X fanout480/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold926/X fanout591/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2 fanout449/X fanout455/X
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/C VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/X sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/A3
+ sky130_fd_sc_hd__nand2_1
XFILLER_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold1141 hold1141/A VGND VGND VPWR VPWR hold1141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1130 hold1130/A VGND VGND VPWR VPWR hold1130/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__and3_2_B
+ m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/B1
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout69_A fanout71/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__xor2_2_A hold674/A hold398/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xhold1174 hold1174/A VGND VGND VPWR VPWR hold1174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1163 hold1163/A VGND VGND VPWR VPWR hold1163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1185 hold1185/A VGND VGND VPWR VPWR hold1185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1152 hold1152/A VGND VGND VPWR VPWR hold1152/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2_X m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout155/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1134/A sky130_fd_sc_hd__dfxtp_1
Xhold1196 hold1196/A VGND VGND VPWR VPWR hold1196/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__or2_2_B fanout485/X hold135/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__mux2_1_A1 fanout427/X
+ m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/B1 m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/A2
+ VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__a22o_2_B2/A2 sky130_fd_sc_hd__mux2_1
XANTENNA_fanout24_X fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout186/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload19 clkload19/A VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__inv_8
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ba_2_A1
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/X VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__o21ba_1
XFILLER_6_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_11_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold946/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold885/A fanout24/X fanout52/X hold1025/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout256/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1036 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold827/X fanout222/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and2_2_B fanout439/X hold64/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_48_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A0 hold258/A m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout509/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold608/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__xor2_2_A hold1138/A hold344/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_35_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2
+ fanout255/X m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ fanout368/X fanout177/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2/X
+ sky130_fd_sc_hd__a221o_1
Xfanout206 fanout207/X VGND VGND VPWR VPWR fanout206/X sky130_fd_sc_hd__buf_4
Xfanout228 fanout228/A VGND VGND VPWR VPWR fanout228/X sky130_fd_sc_hd__buf_4
Xfanout217 fanout218/X VGND VGND VPWR VPWR fanout217/X sky130_fd_sc_hd__buf_4
Xfanout239 fanout239/A VGND VGND VPWR VPWR fanout239/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout273_A fanout273/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold921/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout538_A fanout539/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout159_X fanout159/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2_A1 m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout440_A fanout441/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_65_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold153/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_1098 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout60/X
+ fanout69/X hold1073/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_50_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout108/X
+ fanout132/X hold1026/A m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold104/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout595/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold271 hold271/A VGND VGND VPWR VPWR hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold260 hold260/A VGND VGND VPWR VPWR hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A VGND VGND VPWR VPWR hold293/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A VGND VGND VPWR VPWR hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout284/X m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout289/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A1_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout189/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__or2_2_A hold434/A fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_45_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold155/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_4_1439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout111/A sky130_fd_sc_hd__and4_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout213/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout402/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1 hold685/A fanout382/X
+ fanout194/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/B1
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout468/X fanout474/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2/B1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0 hold1034/X m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold766/X hold698/X fanout601/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__xnor2_2_A hold375/A hold710/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_6_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A hold985/X
+ VGND VGND VPWR VPWR hold984/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_71_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_1328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A1_S fanout411/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold237/A sky130_fd_sc_hd__dfxtp_1
Xinput6 ui_in[3] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C fanout446/X m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C/B
+ m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C/C VGND VGND VPWR VPWR
+ m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/B sky130_fd_sc_hd__and3_1
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold208/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_block_data.data_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y
+ m_io.data_v_early_sky130_fd_sc_hd__and3_2_C/X m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.data_v_early_sky130_fd_sc_hd__a21oi_2_A2/Y VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor3_1
Xm_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
XFILLER_18_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout194/X m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[14\]\[22\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout176/X fanout272/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout119_A fanout119/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B_A fanout489/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/A m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__xnor2_2_A hold1017/A hold963/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_47_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout279/X m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ fanout350/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_fanout488_A fanout489/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold246/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1029 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[8\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold790/A hold589/X fanout603/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_A_sky130_fd_sc_hd__o211a_2_X
+ fanout451/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1/A2
+ fanout401/X fanout468/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout443_X fanout443/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__xnor2_2_A hold402/A m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_51_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout229/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A1_S fanout323/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A0_S fanout509/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__and2_2_A/B fanout425/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XFILLER_26_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold465/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_26_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout592 fanout594/X VGND VGND VPWR VPWR fanout592/X sky130_fd_sc_hd__buf_2
Xfanout581 fanout582/X VGND VGND VPWR VPWR fanout581/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout570 fanout571/X VGND VGND VPWR VPWR fanout570/X sky130_fd_sc_hd__clkbuf_2
XFILLER_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold205/X fanout335/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__nand2_2_B fanout428/X hold177/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_A_N
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.cmd\[2\]_sky130_fd_sc_hd__nor2_2_A block_last_sky130_fd_sc_hd__a32o_2_B2/A1
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A2 VGND VGND VPWR VPWR m_io.cmd\[2\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/B fanout357/X fanout269/A
+ m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold551/X hold513/X fanout545/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A0 hold156/A m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__a31o_2_A3 fanout447/X fanout480/X
+ hold127/A fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A0 hold75/A m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout502/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_11 ANTENNA_11/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_next\[0\]_sky130_fd_sc_hd__and3_2_B_X fanout303/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A fanout236/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__or2_2_A hold519/A fanout373/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_53_1371 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/B
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
XANTENNA_fanout403_A fanout406/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1103/A hold952/X fanout586/X VGND VGND VPWR VPWR hold953/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/A
+ sky130_fd_sc_hd__inv_2
XFILLER_14_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_S fanout214/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1252/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1/X m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B fanout499/X m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1097/X hold530/X fanout598/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout51_A fanout51/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y fanout272/X m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_800 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_50_clk clkload2/A VGND VGND VPWR VPWR clkload21/A sky130_fd_sc_hd__clkbuf_8
XFILLER_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B fanout434/X hold126/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_8_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_buffer\[20\].m_y_buf m_blake2.m_hash256.g_buffer\[20\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[20\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X fanout482/X fanout611/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X/B1
+ sky130_fd_sc_hd__and3b_1
XANTENNA_m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__and3_2_A_B fanout463/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1255/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XFILLER_79_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_A2
+ fanout377/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/X sky130_fd_sc_hd__xor2_1
XFILLER_59_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_41_clk clkload5/A VGND VGND VPWR VPWR clkbuf_leaf_41_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_33_1208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold804 hold804/A VGND VGND VPWR VPWR hold804/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hash\[1\]_sky130_fd_sc_hd__mux2_1_A1_S fanout430/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1_S fanout203/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold815 hold815/A VGND VGND VPWR VPWR hold815/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 hold837/A VGND VGND VPWR VPWR hold837/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1266/X m_blake2.m_hash256.m_matrix\[8\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout544/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold826 hold826/A VGND VGND VPWR VPWR hold826/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold848 hold848/A VGND VGND VPWR VPWR hold848/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold859 hold859/A VGND VGND VPWR VPWR hold859/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__nand2_2_A_B m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_A_N_sky130_fd_sc_hd__o21ba_2_X
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_4_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold798/X hold582/X fanout584/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__xor2_2_B hold872/A hold357/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
XANTENNA_fanout186_A fanout186/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_700 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout289/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout353_A fanout354/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A fanout621/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout239_X fanout239/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clkload4/A VGND VGND VPWR VPWR clkload31/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout520_A fanout524/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__o22a_2_A1_A2 m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout591/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold633/X m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2
+ fanout283/X m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout288/X fanout354/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout406_X fanout406/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_A1
+ fanout295/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A fanout99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/A fanout609/X input4/X VGND VGND VPWR VPWR m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
XFILLER_0_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B/A
+ hold481/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout54_X fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold692/X m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold944/A fanout110/X fanout150/X hold1251/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold476/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y
+ fanout473/X fanout407/X VGND VGND VPWR VPWR fanout266/A sky130_fd_sc_hd__nand2_4
Xm_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__xnor2_2_A hold1118/A hold428/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_21_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_980 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_clk clkload1/A VGND VGND VPWR VPWR clkbuf_leaf_23_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold405/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__a221o_2_A1 hold595/A fanout275/X
+ m_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__or2_2_A/X fanout185/X fanout271/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ hold990/X VGND VGND VPWR VPWR hold989/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold474/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold689/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_S fanout223/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold496/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__nand2_2_B fanout432/X hold192/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_65_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_Q fanout480/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_1128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout60/X fanout40/X
+ hold574/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[12\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold686/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2 m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A2 m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_clkbuf_leaf_62_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout239/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold738/X fanout226/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold299/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold417/A m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout378/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold881/A fanout58/X fanout34/X m_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_14_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkload13/A sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_44_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[8\]_sky130_fd_sc_hd__or2_2_A_B fanout243/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[3\]_sky130_fd_sc_hd__mux2_1_A0_A0 hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold601 hold601/A VGND VGND VPWR VPWR hold601/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 hold612/A VGND VGND VPWR VPWR hold612/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 hold645/A VGND VGND VPWR VPWR hold645/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold623 hold623/A VGND VGND VPWR VPWR hold623/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout101_A fanout103/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold634 hold634/A VGND VGND VPWR VPWR hold634/X sky130_fd_sc_hd__dlygate4sd3_1
Xblock_last_sky130_fd_sc_hd__a22o_2_B2 fanout463/X block_last_sky130_fd_sc_hd__a22o_2_B2/A2
+ block_last_sky130_fd_sc_hd__a22o_2_B2/B1 hold20/X VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout183/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.v_q\[14\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[14\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold308/A sky130_fd_sc_hd__dfxtp_1
Xhold656 hold656/A VGND VGND VPWR VPWR hold656/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold678 hold678/A VGND VGND VPWR VPWR hold678/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold667 hold667/A VGND VGND VPWR VPWR hold667/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold689 hold689/A VGND VGND VPWR VPWR hold689/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold399/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_15_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ hold812/X VGND VGND VPWR VPWR hold811/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold767/X m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_X fanout189/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A3 m_io.cmd\[5\]_sky130_fd_sc_hd__and2b_2_B/X
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold304/X fanout216/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__a32o_2_A1_B1 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold165/A sky130_fd_sc_hd__dfxtp_1
XFILLER_41_703 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_55_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__nand2_2_A hold858/A fanout349/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_55_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1223/A fanout65/X fanout77/X m_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A0/X
+ m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B/B fanout341/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold1193/A fanout86/X fanout130/X hold1131/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold267/X m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout232/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.v_q\[8\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold837/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/B m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__a22o_2_A1_A2 m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2
+ fanout283/X m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ fanout354/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2/Y
+ sky130_fd_sc_hd__a211oi_1
Xm_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__a21o_2_A1 hold18/X fanout337/X
+ m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
Xm_blake2.m_hash256.v_q\[8\]\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold901/X fanout224/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_659 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout201/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ hold488/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2_A2_N_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ hash\[2\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2/Y m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/A2_N
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout300/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1/A2 m_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold475/A m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout380/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_711 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[2\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold641/X hold571/X fanout605/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold991/X fanout219/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__o21a_2_A1 hold1021/A fanout379/X
+ fanout172/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_80_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A0 hold131/A m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout508/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_1363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold444/X m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_config.ll_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold243/X fanout164/X m_io.m_config.ll_q\[19\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout190/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
XFILLER_9_976 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[13\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold869/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A
+ hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold471/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1219/X fanout206/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1094/X fanout554/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_3_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_3_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold278/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold252/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold807/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold885/X fanout542/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XFILLER_39_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold198/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__mux2_1_A0 hold1077/X m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout28 fanout31/A VGND VGND VPWR VPWR fanout28/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_matrix\[3\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[3\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold491/A sky130_fd_sc_hd__dfxtp_1
Xfanout17 fanout19/A VGND VGND VPWR VPWR fanout17/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold172/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold755/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__xnor2_2_A hold862/A hold583/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xfanout39 fanout39/A VGND VGND VPWR VPWR fanout39/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout149_A fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A hold134/A fanout103/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_2
XFILLER_13_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_4
Xm_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold587/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold59/X fanout335/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout330/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ fanout170/X m_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout251/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[28\]_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_S fanout214/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold420 hold420/A VGND VGND VPWR VPWR hold420/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout407/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold453 hold453/A VGND VGND VPWR VPWR hold453/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[7\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold821/X hold539/X fanout602/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout104_X fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold431 hold431/A VGND VGND VPWR VPWR hold431/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold442 hold442/A VGND VGND VPWR VPWR hold442/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout181/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold475 hold475/A VGND VGND VPWR VPWR hold475/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold464 hold464/A VGND VGND VPWR VPWR hold464/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold486 hold486/A VGND VGND VPWR VPWR hold486/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[5\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold691/X VGND VGND VPWR VPWR hold690/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold1061/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xhold497 hold497/A VGND VGND VPWR VPWR hold497/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A hold217/X
+ VGND VGND VPWR VPWR fanout448/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_3 fanout449/X fanout457/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/C VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_3/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1013/A sky130_fd_sc_hd__dfxtp_1
Xhold1131 hold1131/A VGND VGND VPWR VPWR hold1131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_57_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout473_X fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout158/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1120 hold1120/A VGND VGND VPWR VPWR hold1120/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__or2_2_A hold795/A fanout393/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhold1142 hold1142/A VGND VGND VPWR VPWR hold1142/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout416/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.g_buffer\[21\].m_c_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1164 hold1164/A VGND VGND VPWR VPWR hold1164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1153 hold1153/A VGND VGND VPWR VPWR hold1153/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_2
Xhold1175 hold1175/A VGND VGND VPWR VPWR hold1175/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1197 hold1197/A VGND VGND VPWR VPWR hold1197/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X m_io.m_config.ll_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold334/A sky130_fd_sc_hd__dfxtp_1
Xhold1186 hold1186/A VGND VGND VPWR VPWR hold1186/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A0 hold79/A m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xtt_um_essen_630 VGND VGND VPWR VPWR tt_um_essen_630/HI uio_out[4] sky130_fd_sc_hd__conb_1
XTAP_TAPCELL_ROW_0_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_S fanout234/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout89/X
+ fanout93/X m_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout278/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout410/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1055 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/B m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/D VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold856/A fanout128/X fanout144/X hold1025/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_68_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold549/A fanout60/X fanout72/X hold1079/A m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_23_1004 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold197/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold258/X fanout310/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold328/X m_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout542/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X
+ hold708/A fanout95/X fanout151/X hold522/A m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X/C
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout62/X fanout42/X
+ m_blake2.m_hash256.m_matrix\[14\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_32_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold214/X fanout167/X m_io.m_config.ll_q\[30\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold668/A fanout75/X m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout23/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold1081/A fanout73/X m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__or2_2_B fanout493/X hold105/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and3_2_C fanout446/X fanout478/X
+ hold164/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_A2
+ m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold1049/A fanout125/X fanout89/X hold1071/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__nand2_2_A_B fanout349/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ fanout474/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_A1/Y VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_35_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout207 fanout208/X VGND VGND VPWR VPWR fanout207/X sky130_fd_sc_hd__buf_4
Xfanout229 fanout232/A VGND VGND VPWR VPWR fanout229/X sky130_fd_sc_hd__buf_4
Xfanout218 fanout220/A VGND VGND VPWR VPWR fanout218/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_19_Left_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold46/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_67_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout423/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A0 hold67/A m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout266_A fanout266/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_B
+ m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout271/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout433_A fanout434/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout175/X hold682/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[13\].m_c_buf/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_51_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/A
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/X
+ sky130_fd_sc_hd__or3b_1
XANTENNA_fanout221_X fanout221/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_21_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[13\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1158/A hold1099/X fanout598/X VGND VGND VPWR VPWR hold1159/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold250 hold250/A VGND VGND VPWR VPWR hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B
+ fanout288/A m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xhold261 hold261/A VGND VGND VPWR VPWR hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A VGND VGND VPWR VPWR hold294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A VGND VGND VPWR VPWR hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 hold272/A VGND VGND VPWR VPWR hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold579/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A fanout83/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout165/X m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout621/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ fanout450/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_2
XFILLER_58_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1065/A fanout88/X fanout144/X hold962/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__or2_2_B_A fanout486/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold535/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B fanout491/X m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1/X
+ sky130_fd_sc_hd__a21bo_1
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
Xm_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__xnor2_2_A hold385/A hold809/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A
+ m_blake2.m_hash256.g_buffer\[18\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold339/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__a31o_2_A3 fanout447/X fanout480/X
+ hold202/A fanout520/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_6_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B/X m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_71_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold44/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_68_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 ui_in[4] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XFILLER_37_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__a221o_2_A1 hold1145/A fanout351/X
+ fanout263/X hold514/A fanout269/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_80_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y fanout178/X m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__a21oi_2
XFILLER_40_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[12\]_sky130_fd_sc_hd__or2_2_A hold268/A fanout247/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[12\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1/X m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XFILLER_51_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_60_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__xnor2_2_A hold875/A hold572/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2_sky130_fd_sc_hd__o21bai_2_Y
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ sky130_fd_sc_hd__o21bai_4
Xm_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/A2
+ sky130_fd_sc_hd__o21a_2
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A
+ m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1 fanout445/X m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C/D
+ sky130_fd_sc_hd__and4_1
Xm_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
XFILLER_12_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__inv_2_A m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR hash\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout108/X
+ fanout92/X hold493/A m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold150/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout383_A fanout385/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1
+ fanout418/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR fanout220/A sky130_fd_sc_hd__o21ai_4
XANTENNA_m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[23\].m_c_buf m_blake2.m_hash256.g_buffer\[23\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[23\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_934 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hash\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1 hash\[0\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout61/X
+ fanout39/X m_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_2_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_X fanout269/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold171/X fanout327/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout171_X fanout171/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout550_A fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.res_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.res_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C/B
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_54_1317 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold193/A fanout26/X fanout31/X hold1158/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_875 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_A fanout429/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A_B m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__or2_2_A_B fanout248/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout84_X fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout560 fanout561/X VGND VGND VPWR VPWR fanout560/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout593 fanout594/X VGND VGND VPWR VPWR fanout593/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout582 fanout590/X VGND VGND VPWR VPWR fanout582/X sky130_fd_sc_hd__clkbuf_2
Xfanout571 fanout579/X VGND VGND VPWR VPWR fanout571/X sky130_fd_sc_hd__clkbuf_4
XFILLER_73_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout196/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout19/X hold683/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[11\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout554/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X
+ fanout610/X m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/A2 data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/X
+ m_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold23/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_A2 fanout100/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1251/A fanout591/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold156/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_X m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold1196/A fanout124/X fanout128/X hold1123/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold182/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_A
+ fanout477/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1201/A fanout61/X fanout52/X hold896/A m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout146/X
+ fanout122/X hold11/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_53_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold555/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__o211a_2_C1_B1
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0 hold363/A hash\[1\]_sky130_fd_sc_hd__mux2_1_A1/X
+ fanout363/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold75/X fanout309/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_937 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_767 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_12 ANTENNA_12/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A fanout232/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout131_A fanout131/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A hold1109/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_14_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1_A1 m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold509/X fanout208/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__or2_2_A hold189/A fanout392/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_49_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A0 hold22/A m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1074/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_56_786 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout44_A fanout47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__or2_2_B_A fanout487/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__a221o_2_B2 hold1163/A fanout343/X fanout304/X
+ hold487/A fanout268/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__a221o_2_B2/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_3_7_0_clk_X clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_19_1223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_856 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.f_finished_q_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X
+ VGND VGND VPWR VPWR fanout539/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1_C1 m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[24\].m_y_buf m_blake2.m_hash256.g_buffer\[24\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[24\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_812 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[1\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold193/X hold397/X fanout605/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__a22o_2_A1 hold707/A fanout295/X
+ fanout283/X hold761/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout184/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold500/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xfanout390 fanout391/X VGND VGND VPWR VPWR fanout390/X sky130_fd_sc_hd__clkbuf_2
XFILLER_19_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold739/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xinput10 ui_in[7] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_42_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold816 hold816/A VGND VGND VPWR VPWR hold816/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold805 hold805/A VGND VGND VPWR VPWR hold805/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold827 hold827/A VGND VGND VPWR VPWR hold827/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_55_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold849 hold849/A VGND VGND VPWR VPWR hold849/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 hold838/A VGND VGND VPWR VPWR hold838/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout190/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_51_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_51_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_49_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout346_A fanout361/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_4
XFILLER_52_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[6\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold992/X hold1007/A fanout600/X VGND VGND VPWR VPWR hold993/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold287/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout134_X fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout18/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout232/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout301_X fanout301/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout215/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold477/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_hash\[7\]_sky130_fd_sc_hd__and2_2_B_A fanout442/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold321/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold640/X fanout219/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1_A2
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_63_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout300/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__or2_2_A hold241/A fanout379/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A0 hold117/A m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold673/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold679/X m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout297/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.m_matrix\[13\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1197/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold517/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold591/X m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout301/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[10\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold994/X hold912/X fanout585/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_c_buf\[10\]_sky130_fd_sc_hd__o22a_2_X hold710/A fanout175/X
+ m_blake2.m_hash256.g_c_buf\[10\]_sky130_fd_sc_hd__o22a_2_X/B1 fanout254/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[10\].m_c_buf/A sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold617/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A2 m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[7\].m_c_buf/A sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B/A fanout217/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XFILLER_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[4\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1078/X hold946/X fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B_A fanout429/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2 fanout510/X hold130/A
+ m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/B1 m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
Xm_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/A m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__or2_1
XFILLER_54_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold431/X m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2_X m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_78_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_39_1407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_907 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold325/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold703/A m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__or2_2_B/X fanout380/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XFILLER_72_1000 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_44_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold417/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ hold602/X VGND VGND VPWR VPWR hold601/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_40_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_S fanout154/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold209/A m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__or2_2_B/X fanout367/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y_Y
+ fanout176/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.v_q\[10\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ fanout274/X m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout255/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ sky130_fd_sc_hd__a2bb2o_1
Xhold602 hold602/A VGND VGND VPWR VPWR hold602/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__or4bb_2_C_N
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/C
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/D
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2/B1
+ sky130_fd_sc_hd__or4bb_1
Xm_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold799/X m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__or2_2_B fanout485/X hold76/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xhold624 hold624/A VGND VGND VPWR VPWR hold624/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold613 hold613/A VGND VGND VPWR VPWR hold613/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold635 hold635/A VGND VGND VPWR VPWR hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 hold679/A VGND VGND VPWR VPWR hold679/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 hold657/A VGND VGND VPWR VPWR hold657/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold668 hold668/A VGND VGND VPWR VPWR hold668/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 hold646/A VGND VGND VPWR VPWR hold646/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold666/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_block_data.data_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_io.m_block_data.data_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout296_A fanout299/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold743/X m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout153/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1169/A fanout30/X fanout40/X m_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout463_A fanout465/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_26_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold52/A m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout530/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[12\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold445/X hold708/X fanout604/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout349_X fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout471/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/B1
+ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout251_X fanout251/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold624/A fanout75/X m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout23/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold324/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1273 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1140/X hold1147/A fanout591/X VGND VGND VPWR VPWR hold1141/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold784/X hold1119/A fanout564/X VGND VGND VPWR VPWR hold785/A sky130_fd_sc_hd__mux2_1
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__or2_2_B fanout489/X hold252/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_8_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold783/X fanout549/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold305/X m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout156/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold454/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[2\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[2\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1096/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ ANTENNA_11/DIODE m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[3\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold881/X hold1149/A fanout596/X VGND VGND VPWR VPWR hold882/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X
+ m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A/B fanout393/X fanout238/X
+ m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__a22oi_2_B2/Y VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X/A1
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout277/X m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout289/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_2
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout182/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold475/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout193/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_80_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold131/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[30\]_sky130_fd_sc_hd__nand2_2_A hold1210/A fanout357/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[30\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_13_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold669/X VGND VGND VPWR VPWR hold668/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[8\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold835/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B fanout492/X m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout129/X
+ fanout137/X hold727/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__xor2_2_B hold447/A hold341/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold759/X fanout221/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X_B2_sky130_fd_sc_hd__o21a_2_X
+ hold973/A fanout374/X fanout176/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X/B2
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold10/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/C
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_33_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold993/X VGND VGND VPWR VPWR hold992/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold309/A m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout392/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout461/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_46_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout18 fanout19/A VGND VGND VPWR VPWR fanout18/X sky130_fd_sc_hd__clkbuf_4
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__a311o_2_A1_A2 fanout355/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout29 fanout31/A VGND VGND VPWR VPWR fanout29/X sky130_fd_sc_hd__buf_2
XFILLER_23_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold380/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold28/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1 hold485/A fanout380/X
+ fanout193/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_S fanout217/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__or2_2_A hold244/A fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold108/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_A1
+ fanout403/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout211_A fanout212/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ hold1124/X VGND VGND VPWR VPWR hold1123/A sky130_fd_sc_hd__dfxtp_1
Xhold410 hold410/A VGND VGND VPWR VPWR hold410/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2 m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ fanout261/X fanout306/X hold643/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_1 hold302/A m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout396/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A fanout314/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold432 hold432/A VGND VGND VPWR VPWR hold432/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 hold454/A VGND VGND VPWR VPWR hold454/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold421 hold421/A VGND VGND VPWR VPWR hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold443 hold443/A VGND VGND VPWR VPWR hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 hold487/A VGND VGND VPWR VPWR hold487/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 hold465/A VGND VGND VPWR VPWR hold465/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold476 hold476/A VGND VGND VPWR VPWR hold476/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_S fanout411/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold498 hold498/A VGND VGND VPWR VPWR hold498/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold173/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout299_X fanout299/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_X
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1132 hold1132/A VGND VGND VPWR VPWR hold1132/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1072/A fanout90/X fanout142/X hold1088/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xhold1121 hold1121/A VGND VGND VPWR VPWR hold1121/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold106/A sky130_fd_sc_hd__dfxtp_1
Xhold1110 hold1110/A VGND VGND VPWR VPWR hold1110/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_13_Left_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold142/X fanout341/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xdata_idx\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X hold6/X VGND VGND VPWR
+ VPWR data_idx\[0\]_sky130_fd_sc_hd__and4_2_B/D sky130_fd_sc_hd__dfxtp_1
Xhold1143 hold1143/A VGND VGND VPWR VPWR hold1143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_829 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1154 hold1154/A VGND VGND VPWR VPWR hold1154/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1176 hold1176/A VGND VGND VPWR VPWR hold1176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1165 hold1165/A VGND VGND VPWR VPWR hold1165/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1187 hold1187/A VGND VGND VPWR VPWR hold1187/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1198 hold1198/A VGND VGND VPWR VPWR hold1198/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_38_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_B m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xtt_um_essen_631 VGND VGND VPWR VPWR tt_um_essen_631/HI uio_out[2] sky130_fd_sc_hd__conb_1
XFILLER_54_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[10\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_blake2.m_hash256.m_matrix\[10\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold331/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold79/X fanout335/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[15\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold840/X hold648/X fanout543/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_759 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout351/X m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__a22o_2_A1/X fanout180/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B_A fanout487/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_925 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1222/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ hold409/A m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_61_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[5\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1085/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ fanout360/X m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X fanout257/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/A
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ sky130_fd_sc_hd__nor3_1
XFILLER_49_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1 m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1/A2 m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_37_807 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A0 hold224/A m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout513/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold289/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A0 hold225/A m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout502/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__o21a_2_A1 hold887/A fanout379/X
+ fanout251/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__o21a_1
XFILLER_17_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout199/X m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout257/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2
+ fanout274/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__and2_2_B fanout434/X hold161/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__xnor2_2_A hold405/A hold787/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_14_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[7\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold662/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_A m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_10_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_29_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X hold852/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[14\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XTAP_TAPCELL_ROW_35_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout196/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout208 fanout208/A VGND VGND VPWR VPWR fanout208/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1
+ fanout301/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR fanout208/A sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_35_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1/X
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/B
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.v_q\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0 m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X/A1
+ fanout221/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout219 fanout220/X VGND VGND VPWR VPWR fanout219/X sky130_fd_sc_hd__buf_4
XFILLER_80_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_954 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold144/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_1198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D_sky130_fd_sc_hd__a22o_2_X_B2 hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D_sky130_fd_sc_hd__a22o_2_X_A1 m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold337/X m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold67/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1
+ fanout269/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout161_A fanout163/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout259_A fanout260/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__a221o_2_A1 hold509/A fanout349/X
+ fanout260/X hold1260/A m_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__and3_2_A/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/X sky130_fd_sc_hd__a221o_1
XFILLER_23_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout426_A fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__xnor2_2_A hold266/A hold1226/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_52_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold524/X m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout414/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and3b_2_C m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B
+ fanout481/X m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A VGND VGND
+ VPWR VPWR fanout416/A sky130_fd_sc_hd__and3b_2
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout214_X fanout214/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__inv_2_Y_A
+ fanout463/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold251 hold251/A VGND VGND VPWR VPWR hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hold240/A VGND VGND VPWR VPWR hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xhold262 hold262/A VGND VGND VPWR VPWR hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A0 hold167/A m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold487/X fanout161/X m_io.m_config.ll_q\[17\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xhold284 hold284/A VGND VGND VPWR VPWR hold284/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 hold273/A VGND VGND VPWR VPWR hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A VGND VGND VPWR VPWR hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold898/A fanout115/X fanout141/X hold947/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold929/A fanout51/X fanout39/X hold749/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B fanout449/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_2
XANTENNA_fanout74_A fanout75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1095/X hold849/X fanout555/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_1325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__xnor2_2_A hold304/A hold973/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_58_464 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_818 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout130/X fanout122/X
+ m_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A1
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A0 hold168/A m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[0\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/B2 hold483/X fanout602/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/X fanout614/X VGND VGND VPWR VPWR
+ m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[11\]_sky130_fd_sc_hd__a221o_2_X_B1 m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ data\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout63/X fanout47/X hold970/A VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A_Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold438/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout193/X m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout185/X fanout271/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__mux2_1_A1_S fanout214/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold227/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold698/A fanout135/X fanout119/X hold1099/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput8 ui_in[5] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_49_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout277/X m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout289/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A fanout164/X m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout617/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_data\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_A2
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[14\]\[3\]_sky130_fd_sc_hd__mux2_1_A0 hold961/X m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold911/A fanout50/X fanout38/X hold638/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.g_buffer\[24\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xor2_2_A_A
+ m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold563/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A0 hold195/A m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout611/X VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_59_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_A_sky130_fd_sc_hd__o21a_2_X
+ fanout455/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or4_2_A/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B/A
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ data\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout60/X fanout80/X hold1152/A m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1260/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[5\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1195/X hold1111/X fanout573/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout376_A fanout377/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__o22a_2_B1
+ m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3/X
+ m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/X fanout363/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_buffer\[27\].m_c_buf m_blake2.m_hash256.g_buffer\[27\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[27\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_2_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout203/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_54_1329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout429_X fanout429/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__or2_2_A hold259/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_hash\[2\]_sky130_fd_sc_hd__mux2_1_A1_S fanout430/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout413/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_3_3_0_clk_X clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o32a_2_X_B2
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout550 fanout608/X VGND VGND VPWR VPWR fanout550/X sky130_fd_sc_hd__buf_2
Xfanout583 fanout585/X VGND VGND VPWR VPWR fanout583/X sky130_fd_sc_hd__clkbuf_4
Xfanout561 fanout608/X VGND VGND VPWR VPWR fanout561/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout572 fanout575/X VGND VGND VPWR VPWR fanout572/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__a211oi_2_A1 hold384/A fanout283/X
+ m_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__a22o_2_A1/X fanout379/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__a211oi_2_A1/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
Xfanout594 fanout595/X VGND VGND VPWR VPWR fanout594/X sky130_fd_sc_hd__clkbuf_2
XFILLER_58_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1008 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/A
+ hold480/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_73_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
XFILLER_74_798 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold386/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_38_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_12_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__o211ai_2_A2
+ m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B/X
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A1
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_31_1104 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[3\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1026/X hold975/X fanout547/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XFILLER_6_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_47_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
XFILLER_6_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[13\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/A
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/C
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/X
+ sky130_fd_sc_hd__or4_1
XFILLER_69_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__and2_2_A_A
+ m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_9_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold502/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_B
+ fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ sky130_fd_sc_hd__a21bo_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B
+ fanout473/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR fanout273/A sky130_fd_sc_hd__nor2_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__or2_2_A hold388/A fanout378/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_80_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_13 ANTENNA_13/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_846 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout124_A fanout127/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_S fanout221/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold31/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_65_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A_B m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout493_A fanout494/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold522/X fanout604/X
+ VGND VGND VPWR VPWR hold523/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold22/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout198/X m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout190/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__and3_2_C fanout447/X fanout480/X
+ hold57/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XFILLER_47_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/A m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X/B
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout409/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[8\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold564/X hold702/A fanout562/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__mux2_1_A0 hold286/A m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout381/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_1251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout37_A fanout39/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__nand2_1
XFILLER_32_1402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B fanout460/X fanout461/X
+ hold1180/A VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B/X
+ sky130_fd_sc_hd__or3_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ hold185/X m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__a21oi_2_B1/Y VGND VGND
+ VPWR VPWR hold186/A sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A0 hold264/A m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XFILLER_65_1233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold365/X m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout236/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold423/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ hold773/X VGND VGND VPWR VPWR hold1264/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_buffer\[28\].m_y_buf m_blake2.m_hash256.g_buffer\[28\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[28\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__xnor2_2_A hold999/A hold677/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout380 fanout382/X VGND VGND VPWR VPWR fanout380/X sky130_fd_sc_hd__clkbuf_4
Xfanout391 fanout398/X VGND VGND VPWR VPWR fanout391/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ sky130_fd_sc_hd__or2_1
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A3 m_io.cmd\[2\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y/B
+ sky130_fd_sc_hd__nand2_1
XFILLER_19_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__o221a_2_X
+ hold997/A fanout370/X fanout240/X m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y
+ fanout270/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/D1
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A_sky130_fd_sc_hd__or2_2_X
+ hold1004/A fanout103/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/A
+ sky130_fd_sc_hd__or2_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/A1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_1_Left_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__a22o_2_A1 hold580/A fanout189/X
+ fanout195/X hold870/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__and3_2_A hold238/A fanout464/X fanout394/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold18/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_C_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A/C
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.m_matrix\[10\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold630/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput11 uio_in[0] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_42_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0/X
+ m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[14\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold828 hold828/A VGND VGND VPWR VPWR hold828/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__and2_2_B_A fanout431/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold806 hold806/A VGND VGND VPWR VPWR hold806/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 hold817/A VGND VGND VPWR VPWR hold817/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1019 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold839 hold839/A VGND VGND VPWR VPWR hold839/X sky130_fd_sc_hd__dlygate4sd3_1
Xblock_first_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X fanout610/X block_first_sky130_fd_sc_hd__a32o_2_B2/X
+ VGND VGND VPWR VPWR block_first_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_55_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout210/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_69_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2
+ fanout404/X m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__a211o_2_A1/X
+ m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2/Y
+ sky130_fd_sc_hd__a22oi_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout303/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold338/A m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout367/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B fanout495/X hold219/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_A1
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout593/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_990 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_960 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout241_A fanout243/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C fanout259/X
+ m_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__a221o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C
+ fanout407/X m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout133/X
+ fanout149/X hold613/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__and2_2_B fanout428/X hold114/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__or2_2_B fanout485/X hold117/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout127_X fanout127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[12\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1231/X m_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout551/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold460/X m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold808/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hash\[7\]_sky130_fd_sc_hd__and2_2_B_B hash\[7\]_sky130_fd_sc_hd__and2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B
+ fanout444/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/B1 VGND VGND
+ VPWR VPWR fanout180/A sky130_fd_sc_hd__or2_2
Xm_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold469/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1065/X
+ fanout543/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold117/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold370/X m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold223/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__and2_2_X
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A3 m_io.cmd\[2\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/B1_N
+ sky130_fd_sc_hd__a21oi_1
XFILLER_24_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold480/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_12_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_12_665 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_S fanout215/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1
+ m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2b_2_B/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1/Y
+ VGND VGND VPWR VPWR fanout156/A sky130_fd_sc_hd__nor2_2
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_A
+ fanout477/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold569/A m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout397/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1030 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__o21a_2_A1 hold1232/A fanout388/X
+ fanout173/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold341/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold81/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A0 hold125/A m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
XFILLER_23_919 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold297/A sky130_fd_sc_hd__dfxtp_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__inv_2_Y
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X/A2
+ sky130_fd_sc_hd__clkinv_2
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold757/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold792/X m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold83/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__or2_2_A hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_50_1332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold992/A fanout51/X fanout55/X hold631/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B_A fanout429/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold603 hold603/A VGND VGND VPWR VPWR hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__nand2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.data_v_early_sky130_fd_sc_hd__inv_2_Y fanout308/X VGND VGND VPWR VPWR data_v_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__inv_2
Xhold614 hold614/A VGND VGND VPWR VPWR hold614/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 hold636/A VGND VGND VPWR VPWR hold636/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold625 hold625/A VGND VGND VPWR VPWR hold625/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold669 hold669/A VGND VGND VPWR VPWR hold669/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 hold647/A VGND VGND VPWR VPWR hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 hold658/A VGND VGND VPWR VPWR hold658/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout18/X hold508/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[17\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout191_A fanout192/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold133/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__mux2_1_A0 hold716/X m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold801/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[3\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold762/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold709/X m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout289_A fanout290/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.nn_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__xnor2_2_A hold661/A hold1034/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__a32o_2_A1_A2 fanout346/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold52/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold610/X fanout204/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_908 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
XFILLER_0_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout522/X m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A1_S fanout314/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__xnor2_2_A_B m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout509_X fanout509/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_X fanout411/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__inv_2_Y
+ uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1 VGND VGND VPWR
+ VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_matrix\[5\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ hold919/X VGND VGND VPWR VPWR hold918/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__a221o_2_A1_B2 fanout186/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.g_buffer\[26\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__o21a_2_A1 hold892/A fanout387/X
+ fanout170/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_8_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_io.m_config.ll_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X m_io.m_config.ll_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1105/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_76_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1 hold808/A fanout347/X
+ fanout260/X m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_62_1225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold145/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_62_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_838 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__a211o_2_A1 hold373/A fanout279/X
+ m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__a22o_2_A1/X fanout399/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_75_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_1_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A0 hold51/A m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout501/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout244/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[3\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A ANTENNA_13/DIODE
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.m_matrix\[0\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[0\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/B2
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X
+ fanout232/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_73_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N/A
+ sky130_fd_sc_hd__nor2_1
XFILLER_12_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XFILLER_67_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_37_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[2\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1178/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout425/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_33_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold943/A fanout84/X fanout93/X m_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold309/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N
+ fanout277/X m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout400/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_78_1232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ hold1003/A fanout132/X m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A1
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A2
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A3
+ fanout103/X m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o32ai_4
Xm_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/A
+ m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_46_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y
+ ANTENNA_2/DIODE m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1038/A fanout133/X fanout145/X hold667/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout19 fanout19/A VGND VGND VPWR VPWR fanout19/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__a311o_2_A1_A3 fanout249/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__a22o_2_A1 hold1221/X fanout329/X
+ m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__a22o_2_A1/B1 fanout521/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_C
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold575/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ fanout330/X m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__nand3_1
XFILLER_50_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[4\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold536/X hold1177/A fanout587/X VGND VGND VPWR VPWR hold537/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1091/X fanout224/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold400 hold400/A VGND VGND VPWR VPWR hold400/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold411 hold411/A VGND VGND VPWR VPWR hold411/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 hold444/A VGND VGND VPWR VPWR hold444/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 hold433/A VGND VGND VPWR VPWR hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 hold422/A VGND VGND VPWR VPWR hold422/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ hold1224/A hold829/A m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D
+ sky130_fd_sc_hd__and4_2
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold455 hold455/A VGND VGND VPWR VPWR hold455/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 hold477/A VGND VGND VPWR VPWR hold477/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout223/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold466 hold466/A VGND VGND VPWR VPWR hold466/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold488 hold488/A VGND VGND VPWR VPWR hold488/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A0 hold98/A m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout528/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__o21a_2_X_A1
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xhold499 hold499/A VGND VGND VPWR VPWR hold499/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input9_A ui_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1100 hold1100/A VGND VGND VPWR VPWR hold1100/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_58_668 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout194_X fanout194/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1133 hold1133/A VGND VGND VPWR VPWR hold1133/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_A1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1111 hold1111/A VGND VGND VPWR VPWR hold1111/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1122 hold1122/A VGND VGND VPWR VPWR hold1122/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_79_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1144 hold1144/A VGND VGND VPWR VPWR hold1144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1166 hold1166/A VGND VGND VPWR VPWR hold1166/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold1155 hold1155/A VGND VGND VPWR VPWR hold1155/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout361_X fanout361/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xhold1177 hold1177/A VGND VGND VPWR VPWR hold1177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1188 hold1188/A VGND VGND VPWR VPWR hold1188/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1199 hold1199/A VGND VGND VPWR VPWR hold1199/X sky130_fd_sc_hd__dlygate4sd3_1
Xtt_um_essen_632 VGND VGND VPWR VPWR tt_um_essen_632/HI uio_out[1] sky130_fd_sc_hd__conb_1
XANTENNA_m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1027/A fanout68/X fanout36/X hold700/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_0_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_1 hold1180/A m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_1/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and2_2_X
+ hold1255/A m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout290/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout286/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A1_S fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X m_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__a32o_2_B2/A3 sky130_fd_sc_hd__dfxtp_2
Xm_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__or2_2_A hold289/A fanout247/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X hold269/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout138/X
+ fanout142/X hold902/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold118/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B_A fanout487/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold645/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_49_657 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B/B sky130_fd_sc_hd__dfxtp_1
XFILLER_7_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold224/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__xor2_2_A hold587/A hold263/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XFILLER_45_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold920/X m_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout542/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1188/A fanout32/X fanout76/X hold407/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold225/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_1140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold839/A fanout87/X fanout111/X m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__a22o_2_A1 hold330/A fanout290/X
+ fanout278/X hold499/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__and2_2_B fanout430/X hold102/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_34_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[7\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold944/X hold1056/A fanout592/X VGND VGND VPWR VPWR hold945/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1153/A fanout58/X fanout26/X m_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/A2
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/A3
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/B1
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/X
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1108/X fanout555/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout209 fanout212/X VGND VGND VPWR VPWR fanout209/X sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_35_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold606/A fanout110/X fanout122/X hold16/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_45_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__and2b_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y_A
+ fanout422/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[16\]_sky130_fd_sc_hd__o22a_2_X hold1203/A fanout175/X
+ m_blake2.m_hash256.g_c_buf\[16\]_sky130_fd_sc_hd__o22a_2_X/B1 fanout254/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[16\].m_c_buf/A sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.m_matrix\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1001/X hold865/X fanout593/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_69_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__a221o_2_A1_B2 fanout185/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout154_A fanout156/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__xnor2_2_A hold417/A hold597/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1076/X m_blake2.m_hash256.m_matrix\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout607/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2
+ fanout289/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout321_A fanout323/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout302/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__xor2_2_B hold429/A hold1139/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__or2_2_A hold617/A fanout366/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_17_1377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout419_A fanout420/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_17_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_21_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout207_X fanout207/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold65/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[7\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1073/X hold923/X fanout566/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__and2_2_B_A fanout430/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold230 hold230/A VGND VGND VPWR VPWR hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A VGND VGND VPWR VPWR hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 hold252/A VGND VGND VPWR VPWR hold252/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold296 hold296/A VGND VGND VPWR VPWR hold296/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold167/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold285 hold285/A VGND VGND VPWR VPWR hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A VGND VGND VPWR VPWR hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A VGND VGND VPWR VPWR hold274/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_B1_sky130_fd_sc_hd__or3_2_X_A
+ fanout407/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X
+ m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1054/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_48_clk_X clkbuf_leaf_48_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[29\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold168/X fanout323/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout144/X
+ fanout148/X hold1040/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_26_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout22_X fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout137/X
+ fanout117/X m_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A hold267/A m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_35_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[23\]_sky130_fd_sc_hd__o311a_2_X_C1 fanout355/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1/A2 m_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XFILLER_6_712 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold718/A fanout139/X fanout151/X hold581/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A0 hold86/A m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_A_sky130_fd_sc_hd__o211a_2_X_B1
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1216/A sky130_fd_sc_hd__dfxtp_1
XFILLER_77_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__xnor2_2_A hold475/A hold664/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xinput9 ui_in[6] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_80_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout268/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ hold1217/A m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/A_N
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__xnor2_2_B hold430/A hold449/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_71_clk clkload0/A VGND VGND VPWR VPWR clkbuf_leaf_71_clk/X sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_64_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[14\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold822/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold120/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout419/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/Y
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout85/X fanout149/X
+ m_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_58_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold195/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__mux2_1_A0 hold339/A hash\[6\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout386/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__o21a_2_A1 hold1138/A fanout370/X
+ fanout250/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xhash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_67_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout271_A fanout273/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout195/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A1_S fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_2_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__or2_2_A hold372/A fanout394/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhash\[5\]_sky130_fd_sc_hd__mux2_1_A1 hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout428/X VGND VGND VPWR VPWR hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_4
XANTENNA_fanout157_X fanout157/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_60_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_62_clk clkload2/A VGND VGND VPWR VPWR clkload22/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A0 hold615/A m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold959/X hold871/X fanout542/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X
+ hold546/A fanout359/X fanout182/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_matrix\[14\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1071/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.g_buffer\[30\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A0 hold253/A m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold439/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_1150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1008/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__or3b_2_X
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X/A2
+ sky130_fd_sc_hd__or3b_1
Xfanout551 fanout553/X VGND VGND VPWR VPWR fanout551/X sky130_fd_sc_hd__clkbuf_4
Xfanout540 fanout542/X VGND VGND VPWR VPWR fanout540/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xfanout584 fanout585/X VGND VGND VPWR VPWR fanout584/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_clkbuf_leaf_13_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout573 fanout574/X VGND VGND VPWR VPWR fanout573/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout562 fanout563/X VGND VGND VPWR VPWR fanout562/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_matrix\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1165/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout595 fanout599/X VGND VGND VPWR VPWR fanout595/X sky130_fd_sc_hd__clkbuf_4
XFILLER_46_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold791/X m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_28_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_991 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_53_clk clkload3/A VGND VGND VPWR VPWR clkbuf_leaf_53_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_15_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout188/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout18/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_B
+ fanout249/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_S fanout232/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold363/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A
+ fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[17\]_sky130_fd_sc_hd__or2_2_A hold364/A fanout241/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[17\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__a221o_2_A1 hold777/A fanout347/X
+ fanout259/X ANTENNA_11/DIODE m_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_29_1056 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_C
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/B2 hold508/X fanout560/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold371/X fanout165/X m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_42_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1021 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold73/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_44_clk clkload3/A VGND VGND VPWR VPWR clkbuf_leaf_44_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_75_1076 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_1054 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_23_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
XFILLER_53_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_A
+ fanout477/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ fanout611/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__and2_2_B fanout429/X hold133/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout117_A fanout119/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2b_2_B_A_N
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_729 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout486_A fanout500/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__a21o_2_A1 m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold401/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A_sky130_fd_sc_hd__inv_2_Y/A
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout274_X fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ fanout252/X m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout171/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[24\]_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ hold715/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XANTENNA_fanout441_X fanout441/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold893/A fanout24/X fanout40/X m_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_A1
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__a311o_2_A1 hold904/A fanout354/X
+ fanout249/X m_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__o21a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[14\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a311o_1
Xclkbuf_leaf_35_clk clkload4/A VGND VGND VPWR VPWR clkload32/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout539_X fanout539/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_B2
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout156/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C fanout455/X fanout459/X
+ fanout461/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_matrix\[11\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold613/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_blake2.m_hash256.v_q\[12\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1048/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1142/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold240/X fanout166/X m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_69_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold264/X fanout341/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[4\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold348/X fanout228/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1217/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout381 fanout382/X VGND VGND VPWR VPWR fanout381/X sky130_fd_sc_hd__clkbuf_4
Xfanout370 fanout371/X VGND VGND VPWR VPWR fanout370/X sky130_fd_sc_hd__clkbuf_4
Xfanout392 fanout398/X VGND VGND VPWR VPWR fanout392/X sky130_fd_sc_hd__buf_2
XFILLER_47_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold572/X m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout297/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__or2_2_A/X fanout612/X VGND VGND VPWR VPWR
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold526/A sky130_fd_sc_hd__dfxtp_1
XFILLER_59_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout195/X m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout187/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold398/X m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clkload1/A VGND VGND VPWR VPWR clkbuf_leaf_26_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_62_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_791 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold963/X fanout227/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput12 uio_in[1] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ fanout239/X m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__a221o_2_A1/X m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X
+ fanout273/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/A sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_42_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xhold807 hold807/A VGND VGND VPWR VPWR hold807/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold818 hold818/A VGND VGND VPWR VPWR hold818/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout182/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_4
Xm_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold372/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout353/X m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
Xhold829 hold829/A VGND VGND VPWR VPWR hold829/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__nor2_2_B_A fanout499/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/A
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/X
+ sky130_fd_sc_hd__o21ba_1
Xm_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold450/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold338/X fanout410/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[3\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold729/X hold1253/A fanout600/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1146/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__mux2_1_A0 hold134/X m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/B2
+ fanout588/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.d_q\[12\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xclkbuf_leaf_17_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkload14/A sky130_fd_sc_hd__clkbuf_8
XFILLER_40_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X
+ fanout115/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout156/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold936/A fanout46/X m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_fanout234_A fanout236/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold510/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/B2 hold1261/A m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_21_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout401_A fanout403/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout446/X m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A/Y hash_v_sky130_fd_sc_hd__a211o_2_X/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout489_X fanout489/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ hold1261/A m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__a22o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/X
+ sky130_fd_sc_hd__and4_1
Xm_blake2.m_hash256.m_matrix\[0\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1162/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold245/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X
+ hold1206/A fanout81/X m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a2111o_1
XFILLER_16_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_909 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_677 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold828/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_B
+ fanout249/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_S fanout410/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold885/X m_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout546/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nor2_2_Y_Y
+ m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_3_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold569/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__or2_2_A hold605/A fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold300/A fanout61/X fanout45/X hold1178/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold833/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y/B m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/B sky130_fd_sc_hd__a21o_1
XFILLER_6_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_688 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a211o_2_X
+ m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/X
+ m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A3
+ sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and3_2_C_A fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold125/X fanout338/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold834/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_blake2.m_hash256.v_q\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1212/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_758 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_972 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_72_1079 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nand2_1
Xhold615 hold615/A VGND VGND VPWR VPWR hold615/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 hold604/A VGND VGND VPWR VPWR hold604/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 hold626/A VGND VGND VPWR VPWR hold626/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 hold659/A VGND VGND VPWR VPWR hold659/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_6_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_6_clk/X sky130_fd_sc_hd__clkbuf_8
Xhold637 hold637/A VGND VGND VPWR VPWR hold637/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold388/A sky130_fd_sc_hd__dfxtp_1
Xhold648 hold648/A VGND VGND VPWR VPWR hold648/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A ANTENNA_12/DIODE
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__or2_2_B fanout500/X hold78/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[14\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.round_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A hold410/X
+ VGND VGND VPWR VPWR fanout453/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold751/A sky130_fd_sc_hd__dfxtp_1
Xblock_last_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A block_last_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__xnor2_2_A hold363/A hold1216/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout237/X m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout415/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A0 hold206/A m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout536/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_buffer\[10\].m_y_buf m_blake2.m_hash256.g_buffer\[10\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[10\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__a32o_2_A1_A3 fanout249/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__mux2_1_A0 hold99/A m_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout519/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_c_buf\[19\]_sky130_fd_sc_hd__o22a_2_X hold901/A fanout175/X
+ m_blake2.m_hash256.g_c_buf\[19\]_sky130_fd_sc_hd__o22a_2_X/B1 fanout254/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[19\].m_c_buf/A sky130_fd_sc_hd__o22a_1
XFILLER_26_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold346/X fanout570/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout140/X
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout422/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ hold1254/X m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout616_A fanout621/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout237_X fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold302/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout404_X fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold44/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_8_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout97_A fanout99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1187/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xor2_1
XFILLER_1_879 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__o21a_2_A1 hold1107/A fanout385/X
+ fanout172/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[5\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ hash\[7\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_76_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D_sky130_fd_sc_hd__a22o_2_X_B2 hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D_sky130_fd_sc_hd__a22o_2_X_A1 m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold810/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A hold842/X
+ VGND VGND VPWR VPWR hold841/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload21/A m_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_5_1164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold609/A fanout83/X fanout43/X hold1186/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__and2_2
XANTENNA_fanout52_X fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold51/X fanout312/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold876/X fanout595/X
+ VGND VGND VPWR VPWR hold877/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A hold854/X
+ VGND VGND VPWR VPWR hold853/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_80_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_750 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[14\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1186/X m_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout587/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold456/X fanout545/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X m_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold487/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A0 hold176/A m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__o21a_2_A1 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A/A
+ fanout364/X fanout250/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_79_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_37_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A0 hold49/A m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_33_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout286/X m_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout293/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/A1
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_47_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2
+ fanout355/X m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/X
+ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_46_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o21a_2_A2
+ fanout456/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/X fanout444/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o21a_2_A2/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_S fanout215/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_11_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold401 hold401/A VGND VGND VPWR VPWR hold401/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout18/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold114/A sky130_fd_sc_hd__dfxtp_1
Xhold445 hold445/A VGND VGND VPWR VPWR hold445/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 hold434/A VGND VGND VPWR VPWR hold434/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 hold412/A VGND VGND VPWR VPWR hold412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 hold423/A VGND VGND VPWR VPWR hold423/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold467 hold467/A VGND VGND VPWR VPWR hold467/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 hold478/A VGND VGND VPWR VPWR hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 hold456/A VGND VGND VPWR VPWR hold456/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold98/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X
+ hold564/A fanout129/X fanout92/X hold1176/A m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a221o_1
Xhold489 hold489/A VGND VGND VPWR VPWR hold489/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B/Y m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1123 hold1123/A VGND VGND VPWR VPWR hold1123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1101 hold1101/A VGND VGND VPWR VPWR hold1101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 hold1112/A VGND VGND VPWR VPWR hold1112/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1167 hold1167/A VGND VGND VPWR VPWR hold1167/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1145 hold1145/A VGND VGND VPWR VPWR hold1145/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1134 hold1134/A VGND VGND VPWR VPWR hold1134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1156 hold1156/A VGND VGND VPWR VPWR hold1156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1189 hold1189/A VGND VGND VPWR VPWR hold1189/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_B2 hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_A1 m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[25\]_sky130_fd_sc_hd__nor2_2_A hold1181/A fanout368/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/C1 sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout293/X m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ fanout356/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ sky130_fd_sc_hd__a211o_1
Xhold1178 hold1178/A VGND VGND VPWR VPWR hold1178/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold361/X fanout548/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xtt_um_essen_633 VGND VGND VPWR VPWR tt_um_essen_633/HI uio_out[0] sky130_fd_sc_hd__conb_1
Xtt_um_essen_622 VGND VGND VPWR VPWR tt_um_essen_622/HI uio_oe[6] sky130_fd_sc_hd__conb_1
XANTENNA_fanout354_X fanout354/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold589/X hold841/A fanout603/X VGND VGND VPWR VPWR hold590/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/B sky130_fd_sc_hd__a21oi_2
Xm_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_9_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold436/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold746/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_73_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold990 hold990/A VGND VGND VPWR VPWR hold990/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A0 hold137/A m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold381/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__xnor2_2_B hold1232/A hold692/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_76_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout400/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_9_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_754 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_772 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_S fanout204/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_39_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout256/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_35_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__or2_2_A hold220/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y fanout273/X m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_45_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__or2_1
XFILLER_45_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold1034/A fanout276/X m_blake2.m_hash256.v_q\[14\]\[7\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout186/X fanout272/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1074 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout275/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1014 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.g_buffer\[29\].m_y_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_4
Xm_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__mux2_1_A0 hold490/X m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_A1 m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout147_A fanout147/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X
+ hold1252/A fanout137/X m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/B2
+ sky130_fd_sc_hd__a2111o_1
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_21_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B fanout483/X hold190/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout314_A fanout342/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1038/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B fanout425/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold220 hold220/A VGND VGND VPWR VPWR hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold242/A VGND VGND VPWR VPWR hold242/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_matrix\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold253 hold253/A VGND VGND VPWR VPWR hold253/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold231 hold231/A VGND VGND VPWR VPWR hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A VGND VGND VPWR VPWR hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A VGND VGND VPWR VPWR hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 hold275/A VGND VGND VPWR VPWR hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1 hold526/A fanout350/X
+ fanout260/X m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/B2 fanout268/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N_B1_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold297 hold297/A VGND VGND VPWR VPWR hold297/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_63_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__xnor2_2_A hold610/A hold560/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_73_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X_C
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__inv_2_A/A
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ hold1161/A m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout422/A VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A/A
+ hold633/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[11\]_sky130_fd_sc_hd__a221o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_S fanout221/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_731 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold70/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold86/X fanout317/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold626/A fanout136/X fanout148/X m_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout260/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_1151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold248/A m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__or2_2_B/X fanout374/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout142/X fanout94/X
+ hold1170/A m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1149/A fanout134/X fanout94/X hold955/A m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_64_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold315/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold971/X fanout224/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_58_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold970/X hold1060/A fanout600/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__xnor2_2_A hold309/A hold383/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold592/X m_blake2.m_hash256.v_q\[7\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_2_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout264_A fanout265/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold91/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__or2_2_B fanout487/X hold65/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout431_A fanout443/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1147/X m_blake2.m_hash256.m_matrix\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout591/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold615/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold582/X hold1269/X fanout584/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold108/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and3b_2_C_X fanout416/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold253/X fanout326/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o32a_2_X_A3
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold626/X hold543/X fanout557/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__mux2_1_A0 hold427/A m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout376/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xfanout530 fanout538/X VGND VGND VPWR VPWR fanout530/X sky130_fd_sc_hd__clkbuf_4
Xfanout541 fanout542/X VGND VGND VPWR VPWR fanout541/X sky130_fd_sc_hd__clkbuf_2
Xfanout574 fanout575/X VGND VGND VPWR VPWR fanout574/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_A_N_A_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout552 fanout553/X VGND VGND VPWR VPWR fanout552/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold937/A fanout132/X fanout148/X m_blake2.m_hash256.m_matrix\[11\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout563 fanout564/X VGND VGND VPWR VPWR fanout563/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_c_buf\[5\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout596 fanout599/X VGND VGND VPWR VPWR fanout596/X sky130_fd_sc_hd__clkbuf_4
Xfanout585 fanout590/X VGND VGND VPWR VPWR fanout585/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_C_sky130_fd_sc_hd__o31a_2_X
+ fanout407/X fanout460/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B/C
+ sky130_fd_sc_hd__o31a_1
XFILLER_4_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_25_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/B2 hold894/X fanout549/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_25_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A0 hold135/A m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold429/X m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__a22o_2_A1 hold385/A fanout190/X
+ fanout198/X hold495/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ hold866/X VGND VGND VPWR VPWR hold865/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A hold713/A VGND VGND VPWR
+ VPWR m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
XFILLER_29_1024 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__or2_2_B fanout485/X hold112/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X hold1091/A fanout174/A
+ m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1 m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/C1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[31\].m_c_buf/A sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout173/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__a22o_2_A1 hold478/A fanout191/X
+ fanout199/X hold1157/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__or2_2_B_A fanout489/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout182/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__and3_2_C fanout470/X fanout475/X
+ hold333/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XFILLER_75_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_62_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/A1
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1_sky130_fd_sc_hd__a21o_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_33_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_Y m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdata\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X data\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout18/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_B
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold973/X m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout212/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold414/A fanout113/X fanout149/X hold1125/A m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout420/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout239/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold425/X VGND VGND VPWR VPWR hold952/A sky130_fd_sc_hd__dfxtp_1
Xdata\[4\]_sky130_fd_sc_hd__mux2_1_A1 data\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold179/X
+ fanout559/X VGND VGND VPWR VPWR data\[4\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold825/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold1151/A fanout86/X fanout134/X hold1153/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[5\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1020/X hold1085/A fanout570/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1021/X fanout219/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout479_A fanout480/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_S fanout212/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout267_X fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[14\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[14\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1097/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_D_sky130_fd_sc_hd__o311a_2_X_B1
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold547/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout434_X fanout434/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__a211o_2_A1 hold452/A fanout277/X
+ m_blake2.m_hash256.v_q\[1\]\[17\]_sky130_fd_sc_hd__a22o_2_A1/X fanout362/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_71_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A/B fanout206/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout307/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[57\]_sky130_fd_sc_hd__o21a_2_A1 hold159/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/X m_blake2.m_hash256.block_idx_plus_one_q\[57\]_sky130_fd_sc_hd__o21a_2_A1/B1
+ VGND VGND VPWR VPWR hold160/A sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout199/X m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout191/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__xnor2_2_B hold1077/A hold499/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold687/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout82_X fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ hold1224/X m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ fanout427/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_6_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__and3_2_A m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout464/X fanout384/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
Xfanout371 fanout399/X VGND VGND VPWR VPWR fanout371/X sky130_fd_sc_hd__clkbuf_4
Xfanout360 fanout361/X VGND VGND VPWR VPWR fanout360/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout382 fanout385/X VGND VGND VPWR VPWR fanout382/X sky130_fd_sc_hd__buf_2
Xfanout393 fanout398/X VGND VGND VPWR VPWR fanout393/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold707/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold333/X m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[13\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1036/X m_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout587/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__a22o_2_B1 fanout408/X hold1137/A
+ m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/A fanout249/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__a22o_2_B1/X sky130_fd_sc_hd__a22o_1
XFILLER_62_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_17_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/A_N
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__o311a_2_A1/X m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and3b_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xinput13 uio_in[2] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.m_matrix\[11\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ hold846/X VGND VGND VPWR VPWR hold845/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_buffer\[13\].m_c_buf m_blake2.m_hash256.g_buffer\[13\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[13\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout48/X fanout76/X
+ hold1266/A m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_42_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold527/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold242/X m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold808 hold808/A VGND VGND VPWR VPWR hold808/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 hold819/A VGND VGND VPWR VPWR hold819/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__a221o_2_A1 hold978/A fanout358/X
+ fanout261/X hold1160/A m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__and3_2_A/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_55_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__inv_2
XFILLER_44_1319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__a211o_2_A1 hold479/A fanout280/X
+ m_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__a22o_2_A1/X fanout389/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold209/X m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold263/X m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_1054 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_74_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold871/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1413 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_53_759 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold561/X m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1 hold1234/A fanout358/X
+ fanout262/X m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/B2 fanout269/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_984 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1176/A fanout80/X fanout64/X hold654/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_60_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout227_A fanout228/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1155/A fanout117/X fanout93/X m_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1113/X
+ fanout548/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_27_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold355/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold887/X m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout156/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[2\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold705/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout370/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_27_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B/A
+ sky130_fd_sc_hd__nor2_2
XTAP_TAPCELL_ROW_27_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D_sky130_fd_sc_hd__a22o_2_X m_io.m_config.data_i\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1
+ hash\[6\]_sky130_fd_sc_hd__or2_2_B/B VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y
+ fanout173/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold291/X fanout165/X m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ fanout239/X m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y/B sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_12_689 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XFILLER_7_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B fanout495/X hold227/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[8\]\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold710/X fanout221/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A0 hold85/A m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X hash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5/D sky130_fd_sc_hd__a21o_1
XFILLER_65_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A/X fanout612/X VGND VGND VPWR VPWR
+ m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2/Y
+ m_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout402/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
Xfanout190 fanout192/A VGND VGND VPWR VPWR fanout190/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_matrix\[6\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold783/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and3_2_C_B fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkload5_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_792 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[8\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ hold408/X VGND VGND VPWR VPWR hold856/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
Xhold605 hold605/A VGND VGND VPWR VPWR hold605/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 hold627/A VGND VGND VPWR VPWR hold627/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold1101/A fanout136/X m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/B1
+ sky130_fd_sc_hd__a2111o_1
Xhold616 hold616/A VGND VGND VPWR VPWR hold616/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold649 hold649/A VGND VGND VPWR VPWR hold649/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 hold638/A VGND VGND VPWR VPWR hold638/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/B
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold746/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold994/A fanout54/X fanout70/X m_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__or2_2_A/A fanout166/X m_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout620/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold206/X fanout340/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__a22o_2_B1_A1 fanout408/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__a22o_2_B1_B2 fanout249/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold861/A fanout118/X fanout150/X m_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout177_A fanout180/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout559/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold99/X fanout326/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout100/X m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o32a_4
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B/X
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XFILLER_0_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_buffer\[14\].m_y_buf m_blake2.m_hash256.g_buffer\[14\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[14\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_1171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_data\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_932 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout612/X VGND VGND VPWR VPWR m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_55_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout132_X fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout511_A fanout539/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout143/X
+ fanout99/X m_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout271/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__xor2_2_A hold982/A hold509/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_5_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__xnor2_2_A hold286/A hold961/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_770 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X m_io.m_config.ll_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold528/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__or2_2_A hold1086/A fanout388/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout415/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1022/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1263/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_A2
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold176/X fanout338/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout249/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold49/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_79_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_33_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__xor2_2_B hold671/A hold570/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__a22o_2_A1 hold561/A fanout295/X
+ fanout283/X hold462/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_840 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_S
+ fanout430/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_A_N
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold757/X hold718/X fanout573/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.g_buffer\[3\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X
+ hold497/A fanout118/X fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a21o_1
Xhold402 hold402/A VGND VGND VPWR VPWR hold402/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout90/X fanout150/X
+ m_blake2.m_hash256.m_matrix\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold424 hold424/A VGND VGND VPWR VPWR hold424/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_S fanout409/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold435 hold435/A VGND VGND VPWR VPWR hold435/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold413 hold413/A VGND VGND VPWR VPWR hold413/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__mux2_1_A0 hold713/A m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout536/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold457 hold457/A VGND VGND VPWR VPWR hold457/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y
+ hold940/A fanout368/X fanout185/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/A1
+ sky130_fd_sc_hd__o21ai_1
Xhold446 hold446/A VGND VGND VPWR VPWR hold446/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold643/A sky130_fd_sc_hd__dfxtp_1
Xhold468 hold468/A VGND VGND VPWR VPWR hold468/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold479 hold479/A VGND VGND VPWR VPWR hold479/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout519/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout294_A fanout295/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1067/A hold847/X fanout594/X VGND VGND VPWR VPWR hold848/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__xnor2_2_A hold338/A hold941/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold1113 hold1113/A VGND VGND VPWR VPWR hold1113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1102 hold1102/A VGND VGND VPWR VPWR hold1102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1124 hold1124/A VGND VGND VPWR VPWR hold1124/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout181/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1135 hold1135/A VGND VGND VPWR VPWR hold1135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1157 hold1157/A VGND VGND VPWR VPWR hold1157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1146 hold1146/A VGND VGND VPWR VPWR hold1146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1168 hold1168/A VGND VGND VPWR VPWR hold1168/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1179 hold1179/A VGND VGND VPWR VPWR hold1179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xtt_um_essen_623 VGND VGND VPWR VPWR tt_um_essen_623/HI uio_oe[5] sky130_fd_sc_hd__conb_1
Xtt_um_essen_634 VGND VGND VPWR VPWR uio_oe[7] tt_um_essen_634/LO sky130_fd_sc_hd__conb_1
XFILLER_54_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__a22oi_2_B2 hold159/A fanout261/X fanout306/X
+ m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ sky130_fd_sc_hd__a22oi_1
Xm_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_53_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_0_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1073 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.res_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X
+ fanout478/X m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.res_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__or2_2_B fanout487/X hold128/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout284/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2 m_blake2.m_hash256.v_q\[9\]\[9\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout250/X m_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__o21a_2_A1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[9\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a32o_2_X
+ fanout463/X m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A/Y hash_v_sky130_fd_sc_hd__a211o_2_X/A2
+ m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A/X
+ fanout478/X VGND VGND VPWR VPWR m_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/A2
+ sky130_fd_sc_hd__a32o_1
XANTENNA_m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__nand2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_S fanout420/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
XFILLER_22_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_795 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout194/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout34/X fanout78/X
+ hold739/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[17\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1012/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_29_1409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[8\]_sky130_fd_sc_hd__or2_2_A hold1257/X fanout243/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[8\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xhold991 hold991/A VGND VGND VPWR VPWR hold991/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold980 hold980/A VGND VGND VPWR VPWR hold980/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold137/X fanout310/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_62_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout88/X fanout92/X
+ hold1231/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__xnor2_2_A hold370/A hold906/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_75_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[11\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout294/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_740 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[16\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A0 hold82/A m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_777 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout292/X m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ fanout356/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__or2_2_A hold275/A fanout395/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_60_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold763/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_39_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__xnor2_2_A hold569/A hold1114/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_35_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A0 hold35/A m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2
+ fanout266/A m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout400/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.v_q\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1092/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout231/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1064 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1057/A fanout58/X fanout70/X hold998/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1251/X hold1256/A fanout591/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__xnor2_2_A hold416/A hold348/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C/B
+ m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/C sky130_fd_sc_hd__a21o_1
XFILLER_52_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[15\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1164/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[4\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1016/X hold943/X fanout568/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_17_Left_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_21_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout307_A fanout307/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hash\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_Q hash\[0\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold210 hold210/A VGND VGND VPWR VPWR hold210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A VGND VGND VPWR VPWR hold243/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/A VGND VGND VPWR VPWR hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 hold232/A VGND VGND VPWR VPWR hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 hold265/A VGND VGND VPWR VPWR hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 hold276/A VGND VGND VPWR VPWR hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 hold254/A VGND VGND VPWR VPWR hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__nand2_2
Xhold287 hold287/A VGND VGND VPWR VPWR hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_59_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold298 hold298/A VGND VGND VPWR VPWR hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_957 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2
+ fanout403/X m_blake2.m_hash256.v_q\[0\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__a211o_2_A1/X
+ m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a22oi_4
XFILLER_63_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__or2_2_A hold487/A fanout241/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_45_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_843 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__and3_2_A_B fanout465/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[23\]_sky130_fd_sc_hd__o311a_2_X_A1 fanout477/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout24/X fanout28/X
+ hold1053/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A0 hold80/A m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_1359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload23/A m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.fsm_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.fsm_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout422/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A hold354/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_75_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[12\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold609/X m_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout587/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N_B
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[9\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold750/X hold667/X fanout575/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold766/A fanout59/X fanout47/X hold641/A m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A2
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
XFILLER_40_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__and3_2_A hold233/A fanout464/X fanout392/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_1226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_S fanout155/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1007/X hold758/X fanout600/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__a221o_2_A1 hold1037/A fanout251/X
+ fanout172/X hold991/A m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[30\]_sky130_fd_sc_hd__a22o_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_15_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X/A1
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_58_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_721 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_754 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__a22o_2_A1 hold1139/A fanout277/X
+ fanout284/X hold740/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ sky130_fd_sc_hd__nor2_1
XFILLER_3_1422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout189/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/A
+ m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/B m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/X sky130_fd_sc_hd__or3_1
XFILLER_24_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout257_A fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1025/X hold962/X fanout540/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout424_A fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR fanout39/A sky130_fd_sc_hd__nor2_2
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1007 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout212_X fanout212/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_70_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold395/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__o211ai_2_A2_C1
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout520 fanout524/X VGND VGND VPWR VPWR fanout520/X sky130_fd_sc_hd__clkbuf_4
Xfanout531 fanout538/X VGND VGND VPWR VPWR fanout531/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout542 fanout546/X VGND VGND VPWR VPWR fanout542/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout575 fanout579/X VGND VGND VPWR VPWR fanout575/X sky130_fd_sc_hd__clkbuf_2
Xfanout553 fanout561/X VGND VGND VPWR VPWR fanout553/X sky130_fd_sc_hd__buf_2
XANTENNA_fanout72_A fanout75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout564 fanout567/X VGND VGND VPWR VPWR fanout564/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/A1
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A1
+ sky130_fd_sc_hd__or3b_1
Xfanout597 fanout599/X VGND VGND VPWR VPWR fanout597/X sky130_fd_sc_hd__clkbuf_2
Xfanout586 fanout589/X VGND VGND VPWR VPWR fanout586/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2
+ fanout290/X m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout278/X hash\[0\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_hash\[4\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_A fanout403/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_982 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1128/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold996/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_952 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout131/X
+ fanout139/X hold641/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1_sky130_fd_sc_hd__a22o_2_X
+ hold957/A fanout132/X fanout96/X m_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y/B1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_25_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold135/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D_sky130_fd_sc_hd__a22o_2_X m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1
+ hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1018/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_12_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1 hold830/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout427/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_35_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__a21o_2_A1 hold105/X fanout327/X
+ m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B fanout489/X m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A_A m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/X
+ hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout314/X VGND VGND VPWR VPWR hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1083/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q data\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout571/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__and2_2_B fanout430/X hold118/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_53_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[8\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ hold1132/X VGND VGND VPWR VPWR hold1131/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1226/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1_B1
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[5\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A/X
+ m_blake2.m_hash256.g_c_buf\[5\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_c_buf\[5\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout175/X hold844/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[5\].m_c_buf/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_79_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout281/X m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout287/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_62_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/A
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_61_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[1\].m_c_buf m_blake2.m_hash256.g_buffer\[1\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[1\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_25_Left_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold1043/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A0 hold47/A m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout534/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1027/A fanout108/X fanout136/X hold1134/A m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold892/X m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhash\[4\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2/Y
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B/Y VGND VGND VPWR
+ VPWR m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/B1
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X
+ hold1165/A fanout124/X m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/B2
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__nand2_2_A hold1135/A fanout351/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[6\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__or2_2_A hold1043/A fanout369/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout405/X m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__a211o_2_A1/X
+ m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A2 sky130_fd_sc_hd__a22o_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold663/X m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout414/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A1_S fanout409/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_34_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__a22o_2_A1 hold426/A fanout191/X
+ fanout199/X hold755/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ fanout239/A m_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout549/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X
+ hold786/A fanout118/X m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y/A
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/A
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout374_A fanout377/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__nand2_2_A hold1148/A fanout353/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[14\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N
+ fanout277/X m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout400/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_28_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[10\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ hold745/X VGND VGND VPWR VPWR hold744/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold221/X m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_993 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_43_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout403/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_838 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout427_X fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B fanout498/X hold176/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X
+ hold393/A fanout347/X fanout181/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__a21o_1
XFILLER_71_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_blake2.m_hash256.g_buffer\[3\].m_y_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold694/X m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout153/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold664/X m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1/B
+ VGND VGND VPWR VPWR fanout67/A sky130_fd_sc_hd__nor2_2
XFILLER_20_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_52_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__o22a_2_A2/B1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ hold316/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1
+ hash\[7\]_sky130_fd_sc_hd__and2_2_B/B VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold472/A m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout380/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold430/X fanout218/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B fanout495/X hold197/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
Xfanout350 fanout361/A VGND VGND VPWR VPWR fanout350/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout383 fanout385/X VGND VGND VPWR VPWR fanout383/X sky130_fd_sc_hd__clkbuf_4
Xfanout361 fanout361/A VGND VGND VPWR VPWR fanout361/X sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_6_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout372 fanout399/X VGND VGND VPWR VPWR fanout372/X sky130_fd_sc_hd__buf_2
Xfanout394 fanout395/X VGND VGND VPWR VPWR fanout394/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold518/X m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X fanout417/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[14\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1072/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_61_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold978/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.m_matrix\[1\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold435/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A/B fanout206/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold580/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__or2_2_X
+ fanout467/X fanout475/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__or2_1
Xinput14 uio_in[4] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
XANTENNA_m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__a22o_2_B2_A2 fanout265/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_70_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold809 hold809/A VGND VGND VPWR VPWR hold809/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1149/X hold1032/A fanout596/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21bai_2_Y
+ m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o21bai_1
XFILLER_7_875 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_buffer\[17\].m_c_buf m_blake2.m_hash256.g_buffer\[17\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[17\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/B2 m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_55_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold874/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout126/X
+ fanout139/X hold970/A m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold949/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold326/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold143/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/B2 hold1264/X fanout578/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold593/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X fanout182/X m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X/A2
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__o21a_1
XFILLER_42_1066 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1026/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X
+ fanout359/X m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X/B1 sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__o22a_2_A2/X
+ hold130/X fanout323/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold824/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3 fanout453/X fanout457/X
+ fanout461/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/X
+ sky130_fd_sc_hd__o41a_1
XFILLER_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout18/X hold459/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[1\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_34_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout404/X m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__a211o_2_A1/X
+ m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A2
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout122_A fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdata\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold239/X fanout308/X VGND VGND VPWR VPWR data\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1056/X m_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout592/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold482/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[5\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[5\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1070/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.g_buffer\[11\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__xnor2_2_A hold339/A hold763/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A0 hold73/A m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout513/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold581/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold571/A fanout138/X fanout142/X hold397/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1/Y m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__mux2_1_A0 hold290/A m_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/A
+ m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1/B2 hold1052/A m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and4_1
XANTENNA_fanout377_X fanout377/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1208/A fanout108/X fanout112/X hold778/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_buffer\[2\].m_y_buf m_blake2.m_hash256.g_buffer\[2\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[2\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_27_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[7\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold566/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A hold1121/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_930 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_S fanout216/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold72/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[9\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1147/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__mux2_1_X
+ hold284/A m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__and2_2_B/X fanout396/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X/A2 sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_4_889 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold85/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout191 fanout192/X VGND VGND VPWR VPWR fanout191/X sky130_fd_sc_hd__buf_2
Xfanout180 fanout180/A VGND VGND VPWR VPWR fanout180/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__a22o_2_A1 hold999/A fanout251/X
+ fanout172/X hold1127/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A/B
+ sky130_fd_sc_hd__nand2b_2
XFILLER_35_716 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__and3_1
XFILLER_15_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold606 hold606/A VGND VGND VPWR VPWR hold606/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 hold617/A VGND VGND VPWR VPWR hold617/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout158/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout18/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold639 hold639/A VGND VGND VPWR VPWR hold639/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold628 hold628/A VGND VGND VPWR VPWR hold628/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A0 hold433/A m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout519/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/Y m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A/B sky130_fd_sc_hd__xor2_1
XFILLER_48_1275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout406/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1000/X hold1002/X fanout569/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_X
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2/Y
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/A
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A_Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ fanout450/X fanout152/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout481/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold939/A fanout41/X fanout37/X hold414/A m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout25/X fanout29/X
+ m_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_1
XFILLER_20_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_922 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_S fanout201/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[18\].m_y_buf m_blake2.m_hash256.g_buffer\[18\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[18\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/B1
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/C
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1 m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__a22o_2_B2/A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout423/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout504_A fanout509/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhash\[0\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C fanout402/X m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y
+ hash\[0\]_sky130_fd_sc_hd__or2_2_B/X VGND VGND VPWR VPWR hash\[0\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_8_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_X fanout494/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold481/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold481/X m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout413/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_57_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/C
+ sky130_fd_sc_hd__nand3_1
XFILLER_5_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2_sky130_fd_sc_hd__nand2_2_Y_Y
+ fanout267/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__or2_2_A hold233/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[55\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold609/A fanout95/X fanout123/X data\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1090/A
+ fanout603/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout112/X
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1/B
+ sky130_fd_sc_hd__nand2b_2
XFILLER_13_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1
+ fanout286/X m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout292/X fanout355/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/B1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/B
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout181/X m_blake2.m_hash256.v_q\[4\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B/Y
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_matrix\[8\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold558/X hold747/A fanout572/X VGND VGND VPWR VPWR hold559/A sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_73_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout86/X fanout142/X
+ hold693/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/B
+ fanout358/X fanout262/X m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ fanout269/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_B
+ m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__nor2_1
Xm_io.m_config.ll_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout163/X m_io.m_config.ll_q\[8\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X VGND
+ VGND VPWR VPWR hold1258/A sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_37_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_682 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0 hold816/X m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout299/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold368/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__and3_2_A m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout463/X fanout373/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_26_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold863/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_S fanout221/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1221/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y fanout271/X m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
Xm_io.m_config.ll_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold1105/X fanout164/X m_io.m_config.ll_q\[11\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X
+ VGND VGND VPWR VPWR hold1106/A sky130_fd_sc_hd__o211a_1
Xhold425 hold425/A VGND VGND VPWR VPWR hold425/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold403 hold403/A VGND VGND VPWR VPWR hold403/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold414 hold414/A VGND VGND VPWR VPWR hold414/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 hold436/A VGND VGND VPWR VPWR hold436/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold469 hold469/A VGND VGND VPWR VPWR hold469/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold447 hold447/A VGND VGND VPWR VPWR hold447/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 hold458/A VGND VGND VPWR VPWR hold458/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.data_v_early_sky130_fd_sc_hd__a21oi_2_A2 hold5/A data_v_sky130_fd_sc_hd__dfxtp_2_Q/D
+ hold1/X VGND VGND VPWR VPWR m_io.data_v_early_sky130_fd_sc_hd__a21oi_2_A2/Y sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__nand2b_2_B_Y fanout361/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1114 hold1114/A VGND VGND VPWR VPWR hold1114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1103 hold1103/A VGND VGND VPWR VPWR hold1103/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a211o_2_X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1/Y m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/C
+ sky130_fd_sc_hd__a211o_1
Xhold1147 hold1147/A VGND VGND VPWR VPWR hold1147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1158 hold1158/A VGND VGND VPWR VPWR hold1158/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout287_A fanout288/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout28/X
+ fanout64/X hold845/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xhold1136 hold1136/A VGND VGND VPWR VPWR hold1136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1125 hold1125/A VGND VGND VPWR VPWR hold1125/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_22_1212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2
+ fanout163/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1169 hold1169/A VGND VGND VPWR VPWR hold1169/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xtt_um_essen_624 VGND VGND VPWR VPWR tt_um_essen_624/HI uio_oe[4] sky130_fd_sc_hd__conb_1
XFILLER_53_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_c_buf\[22\]_sky130_fd_sc_hd__a2111o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtt_um_essen_635 VGND VGND VPWR VPWR uio_oe[3] tt_um_essen_635/LO sky130_fd_sc_hd__conb_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout621_A input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.kk_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1246/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_0_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout194/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout186/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1 hold143/A m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout499/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__xnor2_2_B hold1239/A hold460/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold970 hold970/A VGND VGND VPWR VPWR hold970/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold981 hold981/A VGND VGND VPWR VPWR hold981/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold992 hold992/A VGND VGND VPWR VPWR hold992/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_1239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input15_A uio_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_479 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1169/X fanout559/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold605/X fanout162/X m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__or2_2_A/X fanout614/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_71_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold84/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_752 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__and2_2_B_A fanout441/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[16\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold330/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[14\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1112/X m_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout563/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold82/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_23_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold219/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout273/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold35/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold265/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_36_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N/Y
+ sky130_fd_sc_hd__nand3b_1
Xclkbuf_leaf_74_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkload9/A sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_69_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.fsm_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and4_2_X_B
+ fanout463/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A0 hold53/A m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout523/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X
+ fanout180/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B fanout434/X hold433/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_15_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_A
+ fanout407/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold211 hold211/A VGND VGND VPWR VPWR hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_X
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A1_N
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold200 hold200/A VGND VGND VPWR VPWR hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold244/A VGND VGND VPWR VPWR hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A VGND VGND VPWR VPWR hold233/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout202_A fanout203/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold222 hold222/A VGND VGND VPWR VPWR hold222/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold266 hold266/A VGND VGND VPWR VPWR hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 hold277/A VGND VGND VPWR VPWR hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold255/A VGND VGND VPWR VPWR hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X/X sky130_fd_sc_hd__xor2_1
Xhold299 hold299/A VGND VGND VPWR VPWR hold299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A VGND VGND VPWR VPWR hold288/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__a32o_2_A1_B1 fanout173/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input7_A ui_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout285/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_X fanout192/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__xnor2_2_B hold1182/A hold709/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_27_811 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A_A m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1 hold394/A fanout382/X
+ fanout186/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_65_clk clkload0/A VGND VGND VPWR VPWR clkload10/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X
+ fanout477/X fanout355/X m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ sky130_fd_sc_hd__and3_4
XFILLER_53_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold222/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold948/A fanout62/X fanout70/X hold820/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_42_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout18/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold80/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout192/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A hold719/X
+ VGND VGND VPWR VPWR hold718/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__a22o_2_A1 hold633/A fanout289/X
+ fanout285/X hold321/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_75_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout423/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XFILLER_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N_C
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout287/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/B1
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__a211oi_2_A1/Y m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2/Y
+ m_blake2.m_hash256.v_q\[0\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X fanout404/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_18_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1 hold1207/A fanout343/X
+ fanout259/X m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout349/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A1_N
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A2_N
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_56_clk clkload3/A VGND VGND VPWR VPWR clkbuf_leaf_56_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1_B2 m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__a22o_2_A1 hold982/A fanout189/X
+ fanout196/X hold805/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y hash\[0\]_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_64_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout145/X
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout182/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout182/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_58_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__or2_2_A hold247/A fanout376/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_67_243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout278/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__mux2_1_A1_S fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_B1
+ fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__and2_2_B_A fanout429/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[6\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1209/X m_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout595/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_47_clk clkload4/A VGND VGND VPWR VPWR clkbuf_leaf_47_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_64_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__nand2b_2_B/Y m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C/Y
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ hold1161/X m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XFILLER_24_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_56_1182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1265/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR fanout31/A sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout58/X fanout70/X
+ m_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[4\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XANTENNA_fanout417_A fanout418/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1253/A fanout86/X fanout131/X hold539/A m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1232/X fanout220/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout205_X fanout205/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[30\]_sky130_fd_sc_hd__a221o_2_A1 hold869/A fanout357/X
+ fanout261/X hold830/A m_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__and3_2_A/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[30\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A1
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout532 fanout538/X VGND VGND VPWR VPWR fanout532/X sky130_fd_sc_hd__clkbuf_2
Xfanout521 fanout524/X VGND VGND VPWR VPWR fanout521/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout510 fanout511/X VGND VGND VPWR VPWR fanout510/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout554 fanout555/X VGND VGND VPWR VPWR fanout554/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xfanout565 fanout566/X VGND VGND VPWR VPWR fanout565/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/A2
+ sky130_fd_sc_hd__or3_1
Xfanout543 fanout545/X VGND VGND VPWR VPWR fanout543/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold987/A sky130_fd_sc_hd__dfxtp_1
Xfanout598 fanout599/X VGND VGND VPWR VPWR fanout598/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout587 fanout589/X VGND VGND VPWR VPWR fanout587/X sky130_fd_sc_hd__clkbuf_4
Xfanout576 fanout578/X VGND VGND VPWR VPWR fanout576/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hash\[4\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_B hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk clkload5/A VGND VGND VPWR VPWR clkbuf_leaf_38_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_61_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31oi_2_Y/B1
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold501/X m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X/B
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_25_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__or2_2_A_B fanout248/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout20_X fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_77_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__xnor2_2_B hold716/A hold462/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__xnor2_2_B/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_A1_N
+ fanout190/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/A2
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout195/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold585/A fanout125/X m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold616/X m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold375/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[1\]_sky130_fd_sc_hd__and2b_2_X m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[1\]_sky130_fd_sc_hd__and2b_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[1\]_sky130_fd_sc_hd__and2b_2_X/X sky130_fd_sc_hd__and2b_1
XFILLER_38_939 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout129/X
+ fanout97/X hold1084/A m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold878/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1_A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clkload4/A VGND VGND VPWR VPWR clkload29/A sky130_fd_sc_hd__clkbuf_8
XFILLER_46_961 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold1171/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold241/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout213/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold756/X m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout158/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_677 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[199\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold47/X fanout338/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold282/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__nand2_2_B fanout436/X hold228/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_buffer\[5\].m_c_buf m_blake2.m_hash256.g_buffer\[5\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[5\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout198/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.m_matrix\[2\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold969/X hold1009/A fanout568/X VGND VGND VPWR VPWR hold1010/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold560/X m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout297/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout193/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[13\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1099/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__or2_2_A hold874/A fanout394/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[12\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1145/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold210/A m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1017/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_714 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/B fanout227/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold852/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_747 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_736 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout367_A fanout371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold634/X hold950/A fanout566/X VGND VGND VPWR VPWR hold635/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1178/A fanout137/X fanout97/X m_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_24_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[9\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold841/X hold938/A fanout603/X VGND VGND VPWR VPWR hold842/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__a22o_2_A1 hold1077/A fanout169/X
+ fanout171/X hold949/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[0\]_sky130_fd_sc_hd__a211o_2_X/A2
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_19_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout155_X fanout155/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout426/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
Xm_blake2.m_hash256.m_matrix\[15\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ hold8/X VGND VGND VPWR VPWR data\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__dfxtp_1
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1177/X m_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout559/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout153/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/B
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__mux2_1_A0_S fanout302/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X
+ fanout127/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_2
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B/A
+ VGND VGND VPWR VPWR fanout63/A sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold917/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__a31o_2_A3 fanout473/X fanout477/X
+ hold688/A fanout378/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold402/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1000/A fanout56/X fanout44/X hold969/A m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold472/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xfanout340 fanout341/X VGND VGND VPWR VPWR fanout340/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout384 fanout385/X VGND VGND VPWR VPWR fanout384/X sky130_fd_sc_hd__clkbuf_2
Xfanout373 fanout374/X VGND VGND VPWR VPWR fanout373/X sky130_fd_sc_hd__buf_2
Xfanout351 fanout353/X VGND VGND VPWR VPWR fanout351/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ fanout475/X VGND VGND VPWR VPWR fanout267/A sky130_fd_sc_hd__nand2_4
Xm_blake2.m_hash256.m_matrix\[10\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold631/X hold581/X fanout573/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout362 fanout365/X VGND VGND VPWR VPWR fanout362/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout395 fanout398/X VGND VGND VPWR VPWR fanout395/X sky130_fd_sc_hd__buf_2
XANTENNA_fanout68_X fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold967/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold149/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_35_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_matrix\[6\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1035/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[7\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold662/X hold634/X fanout566/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_17_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__a21o_2_A1 hold215/X fanout327/X
+ m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__a21o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a21o_1
Xm_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/X fanout609/X input7/X VGND VGND VPWR VPWR m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[8\]\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold787/X fanout223/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1041 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput15 uio_in[5] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__and2_2_B fanout433/X hold100/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[14\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold383/X m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout210/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1096 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold584/A m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout395/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1/X m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_78_850 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1078 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout269/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X/B1
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__o31a_2_A1 hold716/A fanout385/X
+ fanout249/X fanout408/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[5\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__o31a_1
XFILLER_19_994 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1 fanout450/A fanout451/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/C fanout444/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1/X sky130_fd_sc_hd__o31a_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_S fanout416/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_647 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y
+ fanout75/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ hold1224/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 fanout240/X hold528/A
+ m_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XFILLER_14_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold175/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__or2_2_B_A fanout487/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk clkload0/A VGND VGND VPWR VPWR clkbuf_leaf_9_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout115_A fanout115/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold109/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold73/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold290/X fanout309/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout484_A fanout486/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_909 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1094 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_1063 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[6\].m_y_buf m_blake2.m_hash256.g_buffer\[6\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[6\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_52_794 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold497/A fanout30/X fanout54/X hold764/A m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_S fanout411/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_A m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ hold701/X VGND VGND VPWR VPWR hold700/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A1
+ m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold798/A fanout114/X fanout138/X m_blake2.m_hash256.m_matrix\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.ll_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X hold1144/X
+ VGND VGND VPWR VPWR hold317/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__xnor2_2_A hold427/A hold490/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A0 hold166/A m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout527/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/A
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_50_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_S fanout212/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout181 fanout184/X VGND VGND VPWR VPWR fanout181/X sky130_fd_sc_hd__buf_4
Xfanout192 fanout192/A VGND VGND VPWR VPWR fanout192/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout170 fanout170/A VGND VGND VPWR VPWR fanout170/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/X m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__or2_1
XFILLER_74_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[13\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1053/X m_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout563/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_B1
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1045/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_44_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[12\]_sky130_fd_sc_hd__a211o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/X
+ m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__o21ai_2_A1/Y fanout268/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y
+ fanout192/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ hold805/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1/A2 m_blake2.m_hash256.block_idx_plus_one_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xhold607 hold607/A VGND VGND VPWR VPWR hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold187/A sky130_fd_sc_hd__dfxtp_1
Xhold618 hold618/A VGND VGND VPWR VPWR hold618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 hold629/A VGND VGND VPWR VPWR hold629/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[9\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ hold785/X VGND VGND VPWR VPWR hold784/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_1
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold873/A fanout136/X m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__and3_2_C_A fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold416/X m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold29/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_B_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_48_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold433/X fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X
+ fanout248/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.g_buffer\[8\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold330/X m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X fanout300/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1 m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ sky130_fd_sc_hd__nand2_8
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A fanout471/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout232_A fanout232/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X m_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1235/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__o21a_2_A1 hold674/A fanout386/X
+ fanout251/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__o21a_1
XFILLER_18_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_block_last_sky130_fd_sc_hd__a22o_2_B2_A1 fanout463/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2
+ fanout274/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout118_X fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold865/X hold902/A fanout592/X VGND VGND VPWR VPWR hold866/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/C
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A0 hold288/A m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XANTENNA_fanout487_X fanout487/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout299/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and3_2_C_A
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1051 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/Y m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A/B sky130_fd_sc_hd__xnor2_1
XFILLER_5_1112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A_Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold111/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1118/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ sky130_fd_sc_hd__and3_1
XFILLER_10_1375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ sky130_fd_sc_hd__and3_2
XTAP_TAPCELL_ROW_37_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__a22o_2_A1_A2_sky130_fd_sc_hd__and2_2_X_A
+ fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold583/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_33_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__and3_2_A_B fanout465/A VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.g_buffer\[14\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold329/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_62_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_31_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_797 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A0 hold280/A m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout511/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__or2_2_A hold359/A fanout241/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__xnor2_2_A hold242/A hold1023/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold516/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B fanout484/X hold25/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xhold404 hold404/A VGND VGND VPWR VPWR hold404/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 hold426/A VGND VGND VPWR VPWR hold426/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout359/X m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ fanout179/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a211o_1
Xhold415 hold415/A VGND VGND VPWR VPWR hold415/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 hold437/A VGND VGND VPWR VPWR hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 hold459/A VGND VGND VPWR VPWR hold459/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 hold448/A VGND VGND VPWR VPWR hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[5\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold794/X hold690/X fanout585/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1104 hold1104/A VGND VGND VPWR VPWR hold1104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 hold1115/A VGND VGND VPWR VPWR hold1115/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__xnor2_2_A hold209/A hold1018/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold1148 hold1148/A VGND VGND VPWR VPWR hold1148/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1126 hold1126/A VGND VGND VPWR VPWR hold1126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1137 hold1137/A VGND VGND VPWR VPWR hold1137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1159 hold1159/A VGND VGND VPWR VPWR hold1159/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout182_A fanout183/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ hold868/X VGND VGND VPWR VPWR hold867/A sky130_fd_sc_hd__dfxtp_1
Xtt_um_essen_625 VGND VGND VPWR VPWR tt_um_essen_625/HI uio_oe[2] sky130_fd_sc_hd__conb_1
Xm_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__xnor2_2_A hold824/A hold534/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout268/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout447_A fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_S fanout155/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_1017 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout614_A fanout615/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout32/X fanout44/X
+ m_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout235_X fanout235/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/A1
+ m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/A2 m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/Y sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout402_X fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout17/X m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[7\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__xnor2_2_A hold887/A hold489/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_73_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold982 hold982/A VGND VGND VPWR VPWR hold982/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold960 hold960/A VGND VGND VPWR VPWR hold960/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold971 hold971/A VGND VGND VPWR VPWR hold971/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout117/X
+ fanout93/X m_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_915 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold993 hold993/A VGND VGND VPWR VPWR hold993/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout481/X fanout152/X m_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1/B1 m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[113\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_17_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[0\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/A
+ sky130_fd_sc_hd__and2b_1
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_713 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.round_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold409/X fanout152/A m_blake2.m_hash256.round_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ hold1075/A VGND VGND VPWR VPWR hold410/A sky130_fd_sc_hd__o211a_1
XFILLER_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold937/A fanout56/X fanout28/X m_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X
+ fanout359/X m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__a22o_2_A1/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_39_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_A_N m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[12\]_sky130_fd_sc_hd__and2b_2_A_N/X sky130_fd_sc_hd__and2b_1
XANTENNA_m_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__dfxtp_2_Q_Q fanout500/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_985 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_963 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout201/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold938/A fanout34/X fanout43/X m_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold779/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A
+ m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X/B
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/X VGND VGND VPWR VPWR fanout168/A
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_69_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1 m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/B2
+ fanout101/X m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/Y sky130_fd_sc_hd__o22ai_4
Xm_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout568/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold105/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold736/A fanout113/X fanout133/X hold491/A m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold955/A fanout82/X fanout66/X hold1251/A m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_c_buf\[17\]_sky130_fd_sc_hd__a2111o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ fanout459/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
XFILLER_56_1397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold53/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout396/X m_blake2.m_hash256.h_flat\[223\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ m_blake2.m_hash256.v_q\[5\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_1/X fanout191/X fanout179/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__mux2_1_A1_S fanout335/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold201 hold201/A VGND VGND VPWR VPWR hold201/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold238/X fanout166/X m_io.m_config.ll_q\[29\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold862/A sky130_fd_sc_hd__dfxtp_1
Xhold223 hold223/A VGND VGND VPWR VPWR hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A VGND VGND VPWR VPWR hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/A VGND VGND VPWR VPWR hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hold278/A VGND VGND VPWR VPWR hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold245/A VGND VGND VPWR VPWR hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A VGND VGND VPWR VPWR hold256/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold267 hold267/A VGND VGND VPWR VPWR hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold289 hold289/A VGND VGND VPWR VPWR hold289/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[8\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold995/X hold983/X fanout574/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ fanout360/X m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X fanout257/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout397_A fanout398/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout185_X fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__o22a_2_A1 m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2 fanout172/X fanout253/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__o22a_1
XFILLER_22_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_C1 m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_823 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[17\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold809/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold334/X
+ fanout167/X m_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_72_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1225/X fanout207/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold346/A fanout96/X fanout149/X m_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_10_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_c_buf\[23\]_sky130_fd_sc_hd__o311a_2_X_A3 m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[30\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_79_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_S fanout410/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/D
+ fanout422/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_clkbuf_leaf_10_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_75_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_68_1235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xblock_last_sky130_fd_sc_hd__a32o_2_B2 block_last_sky130_fd_sc_hd__a32o_2_B2/A1 block_last_sky130_fd_sc_hd__a32o_2_B2/A2
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A3 block_last_sky130_fd_sc_hd__a32o_2_B2/B1
+ hold20/A VGND VGND VPWR VPWR block_last_sky130_fd_sc_hd__a32o_2_B2/X sky130_fd_sc_hd__a32o_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout577/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold790 hold790/A VGND VGND VPWR VPWR hold790/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ fanout257/X m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/B1
+ fanout396/X fanout179/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_2_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold170/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout157/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X
+ hold672/A fanout374/X fanout185/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/A
+ sky130_fd_sc_hd__o21a_1
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C_D
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and2_2_B_A fanout430/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[13\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[13\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1155/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__xor2_2_A hold593/A hold679/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold165/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout411/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__a22o_2_A1 hold591/A fanout291/X
+ fanout285/X hold341/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__or2_2_B_X fanout422/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_A1
+ fanout354/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold345/A m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout362/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ hold857/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_68_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1002/A fanout57/X fanout81/X m_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout550/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A0 hold103/A m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout521/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_A
+ fanout615/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X
+ fanout276/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold1239/X m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout236/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1/B1 m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
XFILLER_3_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold581/X hold503/X fanout574/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold883/A fanout84/X fanout116/X hold1011/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold452/X m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout413/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_51_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout145_A fanout147/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold642/X fanout164/X m_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__or2_2_A/X fanout617/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A_B m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout312_A fanout314/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__a22o_2_A1 hold799/A fanout189/X
+ fanout197/X hold801/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__or2_2_B fanout495/X hold200/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout100_X fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold631/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_70_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__nand2_2_A hold714/A fanout347/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[19\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xfanout500 fanout500/A VGND VGND VPWR VPWR fanout500/X sky130_fd_sc_hd__buf_2
Xfanout522 fanout524/X VGND VGND VPWR VPWR fanout522/X sky130_fd_sc_hd__clkbuf_4
Xfanout533 fanout534/X VGND VGND VPWR VPWR fanout533/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold248/X m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__o31a_2_A2_B1 fanout249/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout511 fanout539/X VGND VGND VPWR VPWR fanout511/X sky130_fd_sc_hd__clkbuf_4
XFILLER_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout555 fanout561/X VGND VGND VPWR VPWR fanout555/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout566 fanout567/X VGND VGND VPWR VPWR fanout566/X sky130_fd_sc_hd__clkbuf_4
Xfanout544 fanout545/X VGND VGND VPWR VPWR fanout544/X sky130_fd_sc_hd__clkbuf_2
Xfanout599 fanout608/X VGND VGND VPWR VPWR fanout599/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout588 fanout589/X VGND VGND VPWR VPWR fanout588/X sky130_fd_sc_hd__clkbuf_4
Xfanout577 fanout578/X VGND VGND VPWR VPWR fanout577/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C
+ ANTENNA_2/DIODE m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A_sky130_fd_sc_hd__inv_2_Y/A
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold489/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_41_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.g_buffer\[8\].m_y_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_27_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N
+ fanout404/X m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__a211oi_2_A1/Y
+ m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N/X
+ sky130_fd_sc_hd__o2bb2a_1
Xm_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold1114/X m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1152/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold447/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold774/A m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout375/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold681/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1100/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1176/X m_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout562/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold56/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold385/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[22\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1181/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_53_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[6\]_sky130_fd_sc_hd__or2_2_B_A fanout500/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold942/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_66_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold478/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[1\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A hold554/X
+ VGND VGND VPWR VPWR hold553/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold473/X m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout301/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_66_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__and2_2_B_A fanout434/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A0_S fanout520/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_S fanout213/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_987 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold872/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold1107/X fanout219/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold595/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A2
+ sky130_fd_sc_hd__nand2_2
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold766/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold875/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_buffer\[9\].m_c_buf m_blake2.m_hash256.g_buffer\[9\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[9\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold147/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold411/X m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ sky130_fd_sc_hd__dfxtp_4
Xm_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold210/X fanout309/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold860/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/B2 sky130_fd_sc_hd__dfxtp_1
XFILLER_37_962 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[11\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[11\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1125/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[13\]\[11\]_sky130_fd_sc_hd__nor2_2_A hold1023/A fanout377/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/C1 sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B fanout486/X m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[129\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_matrix\[5\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ hold899/X VGND VGND VPWR VPWR hold898/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X_C1
+ fanout271/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold548/X m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout160/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout278/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1044/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout148_X fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_11_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.g_buffer\[16\].m_c_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[11\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1251/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__o21a_2_A1 hold576/A fanout372/X
+ fanout169/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[12\]_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A hold426/A m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout18/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_818 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold83/A m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout530/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xfanout330 fanout342/X VGND VGND VPWR VPWR fanout330/X sky130_fd_sc_hd__buf_2
Xfanout341 fanout342/X VGND VGND VPWR VPWR fanout341/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y fanout273/X m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y/B1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[6\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xfanout352 fanout353/X VGND VGND VPWR VPWR fanout352/X sky130_fd_sc_hd__clkbuf_2
Xfanout374 fanout377/X VGND VGND VPWR VPWR fanout374/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1/X
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xfanout363 fanout365/X VGND VGND VPWR VPWR fanout363/X sky130_fd_sc_hd__clkbuf_4
XFILLER_28_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[0\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/B2 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout385 fanout399/X VGND VGND VPWR VPWR fanout385/X sky130_fd_sc_hd__clkbuf_4
Xfanout396 fanout397/X VGND VGND VPWR VPWR fanout396/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout193/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_B1
+ fanout346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/B1
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_B
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold435/A fanout24/X fanout40/X m_blake2.m_hash256.m_matrix\[14\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_S fanout204/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold262/X m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout154/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_42_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_1340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_59_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold584/X fanout214/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhash\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hash\[0\]_sky130_fd_sc_hd__or2_2_B/B fanout309/X VGND VGND VPWR VPWR hash\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_55_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_42_1013 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__or2_2_A hold262/A fanout372/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout48/X fanout44/X
+ hold1101/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[4\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[4\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1016/A sky130_fd_sc_hd__dfxtp_1
XFILLER_53_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout287/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[8\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold827/A sky130_fd_sc_hd__dfxtp_1
XFILLER_80_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[8\]\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold597/X fanout224/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold967/X hold958/X fanout584/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__a221o_2_A1_B2 fanout185/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout127/X fanout119/X
+ m_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_1115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A0 hold138/A m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout501/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_1284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ fanout256/X m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/B1
+ fanout376/X fanout178/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__a21oi_2_B1 m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ hash\[1\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout242/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout108_A fanout111/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1243/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.g_d\[20\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_64_1282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_704 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_726 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold357/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout265_X fanout265/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[8\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold847/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_S fanout224/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout432_X fanout432/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1089/X m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout155/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__and2_2
Xm_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[231\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold153/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold52/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold104/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[31\]_sky130_fd_sc_hd__mux2_1_A1_S fanout228/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold250/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X
+ fanout188/X m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__and2_2_B/X fanout274/X
+ m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__nor2_2_B/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout80_X fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold166/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[9\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold369/X hold764/X fanout583/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_A1 m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__nand2_2_B fanout437/X hold141/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[102\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__or2_2_A hold1150/A fanout369/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xfanout160 fanout160/A VGND VGND VPWR VPWR fanout160/X sky130_fd_sc_hd__buf_4
XFILLER_47_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout182 fanout183/X VGND VGND VPWR VPWR fanout182/X sky130_fd_sc_hd__buf_6
XFILLER_43_1366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout171 fanout173/A VGND VGND VPWR VPWR fanout171/X sky130_fd_sc_hd__clkbuf_4
XFILLER_74_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout193 fanout194/A VGND VGND VPWR VPWR fanout193/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_47_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/A1
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y/B m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_2
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_48_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout577/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_932 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1/B
+ VGND VGND VPWR VPWR fanout200/A sky130_fd_sc_hd__nor2_4
XTAP_TAPCELL_ROW_48_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_902 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_44_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_44_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/X
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_2
XFILLER_15_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_1326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1060/X hold1005/X fanout602/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout221/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold608 hold608/A VGND VGND VPWR VPWR hold608/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[10\]\[6\]_sky130_fd_sc_hd__o21a_2_A1 hold671/A fanout387/X
+ fanout170/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[6\]_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1 m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ fanout451/X fanout250/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold619 hold619/A VGND VGND VPWR VPWR hold619/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1
+ fanout400/X m_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout266/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__and3_2_C_B fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0 hold247/X m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold675/X m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout569/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__xnor2_2_A hold878/A hold726/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_66_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_4_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold880/A fanout124/X fanout112/X hold768/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__or2_2_B_A fanout487/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold208/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__a22oi_2_B2 m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ fanout261/X fanout306/X hold259/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ sky130_fd_sc_hd__a22oi_1
Xm_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1
+ fanout266/X m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout267/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ sky130_fd_sc_hd__o22a_1
Xdata\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold15/X fanout308/X VGND VGND VPWR VPWR data\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold758/X hold520/X fanout600/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_1081 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout195/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold132/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout225_A fanout228/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XFILLER_1_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_8_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout127/X
+ fanout98/X hold911/A m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X/B
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[58\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold288/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__a31o_2_B1 m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B
+ m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2_B1_sky130_fd_sc_hd__nand2_2_Y_Y
+ fanout240/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B fanout487/X hold19/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_25_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A hold221/A m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_17_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold581/A fanout66/X fanout79/X hold539/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_25_740 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.h_flat\[16\]_sky130_fd_sc_hd__o22a_2_A2/X hold96/X fanout309/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold414/X m_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout572/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X m_io.m_config.ll_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold244/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_49_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A0 hold30/A m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_456 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_2
XFILLER_32_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
XFILLER_32_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout144/X
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout104/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y/A1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_67_1119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__xnor2_2_A hold472/A hold394/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout216/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold11/X fanout593/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_37_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_37_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/D m_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1 hold664/A fanout380/X
+ fanout186/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__xnor2_2_B hold908/A hold333/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout301/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkload3_A clkload3/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold561/A sky130_fd_sc_hd__dfxtp_1
XFILLER_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold205/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_784 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold280/X fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A fanout450/X fanout461/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_2
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold416 hold416/A VGND VGND VPWR VPWR hold416/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold427 hold427/A VGND VGND VPWR VPWR hold427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 hold405/A VGND VGND VPWR VPWR hold405/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 hold449/A VGND VGND VPWR VPWR hold449/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 hold438/A VGND VGND VPWR VPWR hold438/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1105 hold1105/A VGND VGND VPWR VPWR hold1105/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1149 hold1149/A VGND VGND VPWR VPWR hold1149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1138 hold1138/A VGND VGND VPWR VPWR hold1138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1116 hold1116/A VGND VGND VPWR VPWR hold1116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_39_854 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1127 hold1127/A VGND VGND VPWR VPWR hold1127/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_c_buf\[6\]_sky130_fd_sc_hd__a211o_2_X m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__o21a_2_A1/X
+ m_blake2.m_hash256.g_c_buf\[6\]_sky130_fd_sc_hd__a211o_2_X/C1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[6\].m_c_buf/A sky130_fd_sc_hd__a211o_1
XFILLER_66_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout234/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A0 hold102/A m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xtt_um_essen_626 VGND VGND VPWR VPWR tt_um_essen_626/HI uio_oe[1] sky130_fd_sc_hd__conb_1
XFILLER_53_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_D_sky130_fd_sc_hd__o311a_2_X
+ fanout459/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/C
+ fanout401/X fanout468/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B/D
+ sky130_fd_sc_hd__o311a_1
Xm_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold71/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout404/X m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__a211o_2_A1/X
+ m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.g_buffer\[20\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout342_A fanout342/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__a31o_2_A3 fanout447/X fanout480/X
+ hold150/A fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_59_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A0 hold25/A m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout607_A fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout228_X fanout228/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold982/X m_blake2.m_hash256.m_g.b_q\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ fanout158/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_77_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout285/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold972 hold972/A VGND VGND VPWR VPWR hold972/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold961 hold961/A VGND VGND VPWR VPWR hold961/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[11\]_sky130_fd_sc_hd__or2_2_A hold505/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[11\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xhold950 hold950/A VGND VGND VPWR VPWR hold950/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_73_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold994 hold994/A VGND VGND VPWR VPWR hold994/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 hold983/A VGND VGND VPWR VPWR hold983/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A1_S fanout341/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold436/X m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_76_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A_sky130_fd_sc_hd__or2_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B_A fanout435/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/X
+ fanout423/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XFILLER_60_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold914/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X/B1
+ m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2b_1
XFILLER_44_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[11\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold654/X m_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout562/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_53_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_38_1265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_X
+ m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout193/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout359/X m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__nor2_1
XFILLER_60_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/C
+ sky130_fd_sc_hd__and2b_1
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_1105 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout299/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold49/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/A
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1 m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A
+ fanout481/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1/X
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_691 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold456/A fanout52/X fanout68/X hold980/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold830/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_1338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold202 hold202/A VGND VGND VPWR VPWR hold202/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/A VGND VGND VPWR VPWR hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A VGND VGND VPWR VPWR hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold235/A VGND VGND VPWR VPWR hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_c_buf\[22\]_sky130_fd_sc_hd__a2111o_2_X hold819/A fanout174/X
+ m_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__o21a_2_A1/X
+ m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__o21a_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[22\].m_c_buf/A sky130_fd_sc_hd__a2111o_1
Xhold246 hold246/A VGND VGND VPWR VPWR hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A VGND VGND VPWR VPWR hold268/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 hold257/A VGND VGND VPWR VPWR hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C/X
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_2
XFILLER_28_1423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__a32o_2_A1_A2 fanout350/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y_A
+ fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold279 hold279/A VGND VGND VPWR VPWR hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout289/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_1369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_59_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout292_A fanout294/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_61_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1011 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout178_X fanout178/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_846 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_35_890 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__xnor2_2_B hold949/A hold518/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__xnor2_2_B/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[178\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold95/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_10_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A2
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/B1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A1
+ sky130_fd_sc_hd__o311a_2
XFILLER_68_1247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o31a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A/B
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__o31a_2
Xhold780 hold780/A VGND VGND VPWR VPWR hold780/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold791 hold791/A VGND VGND VPWR VPWR hold791/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__mux2_1_A0_A1 hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold557/X m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_1005 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_7_1038 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_4_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_813 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_79_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout268/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[57\]_sky130_fd_sc_hd__a21oi_2_A1_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout51/X fanout75/X
+ hold839/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_44_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__mux2_1_A0_S fanout303/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__nor2_2_B_A fanout499/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[11\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_9_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_15_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_A_N
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_9_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold405/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold345/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1_B1
+ fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1
+ fanout473/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR fanout269/A sky130_fd_sc_hd__or2_4
Xm_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold215/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[3\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1032/X hold924/X fanout596/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1267/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1 hold927/A m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1/A2
+ fanout171/X fanout254/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[1\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__nand2_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__and2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__nand2_2_B_A fanout434/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold103/X fanout329/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1139/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_D_sky130_fd_sc_hd__o311a_2_X_B1
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__nor2_1
XFILLER_56_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A fanout449/X fanout454/X
+ fanout460/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A/X sky130_fd_sc_hd__or4_1
XFILLER_51_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/B2
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout138_A fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold738/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__a22o_2_A1 hold792/A fanout292/X
+ fanout286/X hold751/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold1081/A fanout85/X fanout113/X hold1070/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_30_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout305_A fanout307/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold802/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold906/X fanout228/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold266/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold358/A m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout386/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X
+ m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B fanout358/X fanout269/X
+ m_io.m_config.ll_q\[13\]_sky130_fd_sc_hd__a22o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.round_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ fanout458/X fanout152/X m_blake2.m_hash256.round_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout482/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__o31a_2_A2_A1 fanout408/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout512 fanout516/X VGND VGND VPWR VPWR fanout512/X sky130_fd_sc_hd__clkbuf_4
Xfanout523 fanout524/X VGND VGND VPWR VPWR fanout523/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[0\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/A
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/B
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_1
Xfanout501 fanout502/X VGND VGND VPWR VPWR fanout501/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_1144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout534 fanout537/X VGND VGND VPWR VPWR fanout534/X sky130_fd_sc_hd__buf_2
Xfanout556 fanout561/X VGND VGND VPWR VPWR fanout556/X sky130_fd_sc_hd__clkbuf_2
XFILLER_24_1106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout295_X fanout295/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout545 fanout546/X VGND VGND VPWR VPWR fanout545/X sky130_fd_sc_hd__clkbuf_4
Xfanout589 fanout590/X VGND VGND VPWR VPWR fanout589/X sky130_fd_sc_hd__clkbuf_2
Xfanout578 fanout579/X VGND VGND VPWR VPWR fanout578/X sky130_fd_sc_hd__clkbuf_4
XFILLER_24_1139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout567 fanout579/X VGND VGND VPWR VPWR fanout567/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold823/A sky130_fd_sc_hd__dfxtp_1
XFILLER_73_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__and2_2_B fanout428/X hold92/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X/X sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_1_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_805 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold304/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_698 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold466/X m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold952/A fanout82/X fanout66/X hold732/A m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_871 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold774/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold696/X fanout583/X
+ VGND VGND VPWR VPWR hold697/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A_1_A fanout472/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_A1
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold64/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout193/X m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout176/X fanout273/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_57_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold703/X m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold901/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold797/X fanout164/X m_io.m_config.ll_q\[27\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[6\]_sky130_fd_sc_hd__or2_2_B_B hash\[6\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_790 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_719 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_996 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold991/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold268/X
+ fanout167/X m_io.m_config.ll_q\[4\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X VGND
+ VGND VPWR VPWR hold269/A sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold396/A m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout368/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_d\[19\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout190/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1182/X fanout219/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold449/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_S fanout410/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A_Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_71_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A0 hold451/A m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout521/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y_A
+ fanout520/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[13\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1219/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1093/X hold722/X fanout573/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold426/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_708 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold543/A fanout136/X fanout92/X m_blake2.m_hash256.m_matrix\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_64_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_451 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/B m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout255_A fanout258/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_24_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold198/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout161/X m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout611/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout422_A fanout422/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y
+ fanout236/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout183/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__mux2_1_A0 hold281/X m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_39_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A hold925/X
+ VGND VGND VPWR VPWR hold924/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold587/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__xnor2_2_A hold495/A hold816/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_1228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_1206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_4
XANTENNA_m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout291/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold83/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xfanout320 fanout323/X VGND VGND VPWR VPWR fanout320/X sky130_fd_sc_hd__buf_2
XFILLER_78_329 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold788/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout331 fanout332/X VGND VGND VPWR VPWR fanout331/X sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_21_Left_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout342 fanout342/A VGND VGND VPWR VPWR fanout342/X sky130_fd_sc_hd__buf_4
Xfanout375 fanout376/X VGND VGND VPWR VPWR fanout375/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout70_A fanout71/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout353 fanout354/X VGND VGND VPWR VPWR fanout353/X sky130_fd_sc_hd__buf_2
XFILLER_47_705 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout364 fanout365/X VGND VGND VPWR VPWR fanout364/X sky130_fd_sc_hd__dlymetal6s2s_1
Xm_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1080/X fanout572/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout397 fanout398/X VGND VGND VPWR VPWR fanout397/X sky130_fd_sc_hd__clkbuf_4
Xfanout386 fanout388/X VGND VGND VPWR VPWR fanout386/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[12\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout549/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_55_760 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__or2_2_B fanout488/X hold273/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A hold1249/X
+ VGND VGND VPWR VPWR hold1248/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout202/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[14\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1130/X hold1072/X fanout595/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_42_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1190 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_30_Left_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/B1
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_buffer\[22\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A0 hold58/A m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout537/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold461/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_46_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A0 hold126/A m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_42_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_13_1396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold331/A fanout54/X fanout82/X hold1090/A m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout414/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold607/X VGND VGND VPWR VPWR hold606/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_55_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C_D
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1025 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
XFILLER_55_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold258/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_B1
+ fanout239/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout275/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold1037/X m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout155/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold138/X fanout309/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout70/X fanout78/X
+ hold847/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand2_2_B
+ fanout445/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_A1/Y VGND
+ VGND VPWR VPWR fanout152/A sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout183/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_1261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout198/X m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[166\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout190/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_9_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1179/X m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout596/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_749 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout372_A fanout399/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2
+ hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ sky130_fd_sc_hd__a21bo_1
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1/X m_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X
+ fanout273/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_27_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout160_X fanout160/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout258_X fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A0 hold28/A m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
XFILLER_79_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold744/X m_blake2.m_hash256.m_matrix\[10\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout564/X
+ VGND VGND VPWR VPWR hold745/A sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_50_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_50_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A_Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout409/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout161 fanout163/X VGND VGND VPWR VPWR fanout161/X sky130_fd_sc_hd__clkbuf_4
Xfanout150 fanout151/X VGND VGND VPWR VPWR fanout150/X sky130_fd_sc_hd__clkbuf_4
Xm_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__or2_2_A hold246/A fanout243/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xfanout183 fanout184/X VGND VGND VPWR VPWR fanout183/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B fanout483/X hold158/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xfanout172 fanout173/X VGND VGND VPWR VPWR fanout172/X sky130_fd_sc_hd__clkbuf_4
Xfanout194 fanout194/A VGND VGND VPWR VPWR fanout194/X sky130_fd_sc_hd__buf_2
XFILLER_43_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_A2
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_899 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout154/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold999/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_944 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__and3_2_A hold246/A fanout463/X fanout368/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_48_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ fanout475/X VGND VGND VPWR VPWR fanout283/A sky130_fd_sc_hd__nor2_4
Xm_blake2.m_hash256.m_matrix\[8\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold702/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold390/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_44_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__or4_2_B
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__or4_2_B/X
+ sky130_fd_sc_hd__or4_1
XANTENNA_m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_1447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__and3b_2_X_A_N
+ m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold609 hold609/A VGND VGND VPWR VPWR hold609/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1034/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_1245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__xnor2_2_A hold336/A hold1225/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.g_buffer\[19\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout84/X fanout96/X
+ m_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_59_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__xnor2_2_A hold756/A hold915/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_34_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XFILLER_22_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_2
Xm_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B fanout437/X hold50/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__a221o_2_A1 hold851/A fanout344/X
+ fanout259/X hold829/A fanout268/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout120_A fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__xnor2_2_B hold576/A hold663/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout218_A fanout220/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A1_N
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A2_N
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_49_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__xnor2_2_A hold860/A hold1019/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_66_1378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/X
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XFILLER_75_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_877 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold171/A sky130_fd_sc_hd__dfxtp_1
XFILLER_40_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_774 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A1 m_io.cmd\[5\]_sky130_fd_sc_hd__and2b_2_B/X
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1002 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold30/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C/C
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B fanout490/X hold148/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__a31o_2_B1 m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ hold1161/A m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B
+ m_blake2.m_hash256.v_q\[13\]\[19\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_66_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/A1
+ sky130_fd_sc_hd__nand2_1
XFILLER_16_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold127/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ hold495/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_S fanout412/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_766 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout193/X m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout186/X fanout272/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
XFILLER_15_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold936/X fanout598/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_50_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clkload1/A VGND VGND VPWR VPWR clkbuf_leaf_10_clk/X sky130_fd_sc_hd__clkbuf_8
Xhold406 hold406/A VGND VGND VPWR VPWR hold406/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__xnor2_2_A hold584/A hold275/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold417 hold417/A VGND VGND VPWR VPWR hold417/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 hold439/A VGND VGND VPWR VPWR hold439/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold428 hold428/A VGND VGND VPWR VPWR hold428/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__and3_2_C_A fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__o21ai_2_A1 m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[20\]_sky130_fd_sc_hd__a22o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X hold894/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[21\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
Xhold1106 hold1106/A VGND VGND VPWR VPWR hold1106/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__xnor2_4
XANTENNA_hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1 hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1128 hold1128/A VGND VGND VPWR VPWR hold1128/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold156/A sky130_fd_sc_hd__dfxtp_1
Xhold1117 hold1117/A VGND VGND VPWR VPWR hold1117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_26_1384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1139 hold1139/A VGND VGND VPWR VPWR hold1139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_6_1445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_866 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold102/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xtt_um_essen_627 VGND VGND VPWR VPWR tt_um_essen_627/HI uio_oe[0] sky130_fd_sc_hd__conb_1
XANTENNA_m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_A fanout168/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[4\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout576/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold75/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold661/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N/X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout335_A fanout342/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold25/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_788 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout123_X fanout123/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1264/A hold772/X fanout578/X VGND VGND VPWR VPWR hold773/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout502_A fanout509/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o22ai_2_A1
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__nor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ sky130_fd_sc_hd__o22ai_1
XFILLER_33_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhash\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X hash\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[0\]_sky130_fd_sc_hd__or2_2_B/B sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_77_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold940 hold940/A VGND VGND VPWR VPWR hold940/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold973 hold973/A VGND VGND VPWR VPWR hold973/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 hold962/A VGND VGND VPWR VPWR hold962/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold951 hold951/A VGND VGND VPWR VPWR hold951/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout492_X fanout492/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_73_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhash\[1\]_sky130_fd_sc_hd__mux2_1_A1 hash\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0 hash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout430/X VGND VGND VPWR VPWR hash\[1\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_2
XTAP_TAPCELL_ROW_73_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold509/A sky130_fd_sc_hd__dfxtp_1
Xhold995 hold995/A VGND VGND VPWR VPWR hold995/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 hold984/A VGND VGND VPWR VPWR hold984/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_62_1039 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1218/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_68_clk clkload0/A VGND VGND VPWR VPWR clkbuf_leaf_68_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout587/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_814 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout352/X m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X fanout258/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.m_matrix\[14\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[14\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1082/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout36_X fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_B
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__a32o_2_A1 hold482/A fanout350/X
+ fanout252/X fanout173/A m_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__a32o_2_A1/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_40_596 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X hold597/A fanout174/X
+ m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2 hold1046/A m_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[21\].m_c_buf/A sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_39_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__o21ba_2_A1 hold737/A fanout373/X
+ m_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__a22o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[18\]_sky130_fd_sc_hd__o21ba_2_A1/X
+ sky130_fd_sc_hd__o21ba_1
XFILLER_80_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__or2_2_A hold214/A fanout247/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_59_clk clkload2/A VGND VGND VPWR VPWR clkbuf_leaf_59_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_75_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
XANTENNA_m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout614/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__a22o_2_A1 hold398/A fanout294/X
+ fanout286/X hold527/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_35_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_17_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B fanout426/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XFILLER_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N_sky130_fd_sc_hd__and2b_2_X
+ m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__and2_2_A/B m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold203 hold203/A VGND VGND VPWR VPWR hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_68_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold214 hold214/A VGND VGND VPWR VPWR hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold898/X fanout559/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold225 hold225/A VGND VGND VPWR VPWR hold225/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_A m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold269 hold269/A VGND VGND VPWR VPWR hold269/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 hold247/A VGND VGND VPWR VPWR hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/A VGND VGND VPWR VPWR hold236/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xhold258 hold258/A VGND VGND VPWR VPWR hold258/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B_A fanout494/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__a32o_2_A1_A3 fanout252/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__and3_2_X
+ hold2/A hold6/A m_io.data_v_early_sky130_fd_sc_hd__and3_2_C/X VGND VGND VPWR VPWR
+ m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X
+ hold794/A fanout114/X fanout146/X m_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X/C
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y_B
+ fanout407/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold620/A fanout73/X m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout21/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__a21oi_2_B1/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[2\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
XANTENNA_fanout285_A fanout288/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1 hold162/A fanout101/X
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/B1 m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/X
+ sky130_fd_sc_hd__o22a_2
XPHY_EDGE_ROW_77_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[18\]_sky130_fd_sc_hd__mux2_1_A1_S fanout216/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout240_X fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[8\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_769 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1 m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_2
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[3\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold400/X m_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout572/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_75_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A
+ fanout481/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_2
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold633/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X
+ hold351/A fanout103/X m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A1_N
+ sky130_fd_sc_hd__o22a_2
Xhold781 hold781/A VGND VGND VPWR VPWR hold781/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold770 hold770/A VGND VGND VPWR VPWR hold770/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout223/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__nand2_1
XFILLER_49_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold792 hold792/A VGND VGND VPWR VPWR hold792/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1
+ fanout288/X m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout283/X fanout354/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B
+ m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y/B
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ sky130_fd_sc_hd__or3_4
Xm_blake2.m_hash256.m_matrix\[13\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold876/X hold861/X fanout595/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_950 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1/B
+ VGND VGND VPWR VPWR fanout79/A sky130_fd_sc_hd__nor2_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[108\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_18_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[11\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold640/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_825 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input13_A uio_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A hold650/X
+ VGND VGND VPWR VPWR hold649/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_17_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold692/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N_sky130_fd_sc_hd__nor2_2_Y_A
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout417/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout81/X fanout45/X
+ hold1252/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X_C
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y
+ fanout200/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[0\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold907/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold982/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold380/X m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__a22o_2_A1_B2 fanout249/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold534/X m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[13\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1169/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold367/X m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout111/X
+ fanout115/X hold749/A m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/B1 m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D/C
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold770/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B/A sky130_fd_sc_hd__dfxtp_1
XFILLER_55_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_A1_N
+ fanout192/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_S fanout201/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold841/A fanout127/X fanout114/X m_blake2.m_hash256.m_matrix\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[15\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[15\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold720/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2 fanout517/X hold207/A
+ m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/B1 m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__or2_2_B fanout486/X hold132/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1090/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold611/X m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__xor2_2_B hold470/A hold373/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_A_N m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[28\]_sky130_fd_sc_hd__and2b_2_A_N/X sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/A2
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold417/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout271/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout200_A fanout200/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold358/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_70_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1200/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1
+ fanout477/X fanout249/X VGND VGND VPWR VPWR fanout170/A sky130_fd_sc_hd__nor2_1
Xfanout513 fanout516/X VGND VGND VPWR VPWR fanout513/X sky130_fd_sc_hd__buf_2
XFILLER_63_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout524 fanout539/X VGND VGND VPWR VPWR fanout524/X sky130_fd_sc_hd__buf_2
Xfanout502 fanout509/X VGND VGND VPWR VPWR fanout502/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_input5_A ui_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout535 fanout537/X VGND VGND VPWR VPWR fanout535/X sky130_fd_sc_hd__clkbuf_4
XFILLER_63_1167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout557 fanout561/X VGND VGND VPWR VPWR fanout557/X sky130_fd_sc_hd__clkbuf_4
Xfanout546 fanout608/X VGND VGND VPWR VPWR fanout546/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold440/X m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout158/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_63_1189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__a31o_2_B1_A1
+ m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout190_X fanout190/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout579 fanout608/X VGND VGND VPWR VPWR fanout579/X sky130_fd_sc_hd__buf_2
Xfanout568 fanout569/X VGND VGND VPWR VPWR fanout568/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout288_X fanout288/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold767/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_1_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout295/X m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__o21a_2_A1 hold1110/A fanout365/X
+ fanout169/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_io.m_block_data.data_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_io.m_block_data.data_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold6/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout287/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_647 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_989 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_978 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2
+ fanout287/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_883 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout300/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A_1_B fanout407/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold600/A m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout510/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.cmd\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X fanout1/X fanout609/X
+ input13/X VGND VGND VPWR VPWR m_io.cmd\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X hold1055/A fanout276/X m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/C1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/X
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.m_matrix\[0\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[0\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold351/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold267/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_57_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold469/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_1_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0 hold96/A m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout502/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__a31o_2_B1_A3
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_66_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_66_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold674/X m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout155/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold571/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold475/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold396/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__and3_2_A hold218/A fanout464/X fanout395/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[44\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold131/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold451/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xdata_idx\[3\]_sky130_fd_sc_hd__and4_2_A data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/A
+ data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/B data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/C
+ data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/D VGND VGND VPWR VPWR data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/X
+ sky130_fd_sc_hd__and4_1
Xm_blake2.m_hash256.m_matrix\[14\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1082/X m_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout604/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_1421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ hold537/X VGND VGND VPWR VPWR hold536/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold232/X m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout232/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold759/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload20/A m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[8\]\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold941/X fanout221/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[14\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold939/X m_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout572/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A_1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D/C
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__o21ai_2_A1 hold516/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout425/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XFILLER_36_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A2
+ sky130_fd_sc_hd__o31a_2
XANTENNA_fanout150_A fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1147/A fanout34/X fanout66/X hold1256/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/B m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_19_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_A fanout248/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X
+ m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1077/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[6\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1051/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_blake2.m_hash256.round_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout460/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout415_A fanout416/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout203_X fanout203/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold340/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold762/A fanout56/X fanout28/X hold1250/A m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xfanout321 fanout323/X VGND VGND VPWR VPWR fanout321/X sky130_fd_sc_hd__clkbuf_4
XFILLER_8_1123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout332 fanout342/X VGND VGND VPWR VPWR fanout332/X sky130_fd_sc_hd__clkbuf_4
Xfanout310 fanout314/X VGND VGND VPWR VPWR fanout310/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xfanout343 fanout344/X VGND VGND VPWR VPWR fanout343/X sky130_fd_sc_hd__clkbuf_4
Xfanout354 fanout361/A VGND VGND VPWR VPWR fanout354/X sky130_fd_sc_hd__clkbuf_4
Xfanout365 fanout371/X VGND VGND VPWR VPWR fanout365/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_6_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout398 fanout399/X VGND VGND VPWR VPWR fanout398/X sky130_fd_sc_hd__clkbuf_2
Xfanout376 fanout377/X VGND VGND VPWR VPWR fanout376/X sky130_fd_sc_hd__buf_2
Xfanout387 fanout388/X VGND VGND VPWR VPWR fanout387/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 hash\[7\]_sky130_fd_sc_hd__and2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A1 m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__inv_2_A_Y fanout408/A VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold142/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_997 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_27_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X
+ fanout349/X m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__a22o_2_A1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold79/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_C1
+ fanout354/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdata_idx\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X hold2/X VGND VGND VPWR
+ VPWR data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[245\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold58/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_46_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[124\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold126/X fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold424/A fanout94/X fanout122/X hold14/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_42_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[3\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[3\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1002/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__nand2_2_B_A fanout429/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout196/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[5\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold974/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ fanout461/A fanout152/X m_blake2.m_hash256.round_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ fanout482/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[190\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold902/X hold1088/A fanout591/X VGND VGND VPWR VPWR hold903/A sky130_fd_sc_hd__mux2_1
XFILLER_34_901 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
XFILLER_19_953 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__and2_2_B fanout436/X hold921/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_34_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[5\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold414/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__and2_2
XTAP_TAPCELL_ROW_16_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1/Y
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_4
XFILLER_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A0 hold741/A m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout521/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X m_io.m_config.ll_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold291/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A0 hold212/A m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__xnor2_2_A hold345/A hold1203/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__a22o_2_A1 hold879/A fanout174/A
+ m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__or2_2_A/X fanout252/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/B1 sky130_fd_sc_hd__a22o_1
Xm_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout242/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout198_A fanout200/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1/B
+ VGND VGND VPWR VPWR fanout35/A sky130_fd_sc_hd__nor2_2
XFILLER_29_717 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout282/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout18/X m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[24\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XFILLER_37_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout365_A fanout371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold359/X fanout161/X m_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_fanout532_A fanout538/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout153_X fanout153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X m_blake2.m_hash256.h_flat\[54\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold67/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_1380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout418_X fanout418/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold28/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B
+ fanout277/X m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__or2_2_B/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_20_672 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold317/X
+ fanout162/X m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[0\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.m_matrix\[6\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1033/X hold1200/A fanout555/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold897/A fanout141/X fanout120/X m_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__xnor2_2_A hold248/A hold636/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_78_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/A
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ sky130_fd_sc_hd__nor3_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout140 fanout143/X VGND VGND VPWR VPWR fanout140/X sky130_fd_sc_hd__buf_4
Xfanout162 fanout163/X VGND VGND VPWR VPWR fanout162/X sky130_fd_sc_hd__clkbuf_4
Xfanout151 fanout151/A VGND VGND VPWR VPWR fanout151/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout173 fanout173/A VGND VGND VPWR VPWR fanout173/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout195 fanout197/X VGND VGND VPWR VPWR fanout195/X sky130_fd_sc_hd__clkbuf_4
Xfanout184 fanout184/A VGND VGND VPWR VPWR fanout184/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout66_X fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold499/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold220/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A0 hold26/A m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout523/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_70_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout84/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_989 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__xnor2_2_A hold774/A hold389/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A0 hold152/A m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout183/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdata_idx\[0\]_sky130_fd_sc_hd__and4_2_B fanout599/X data_idx\[0\]_sky130_fd_sc_hd__and4_2_B/B
+ data_idx\[0\]_sky130_fd_sc_hd__and4_2_B/C data_idx\[0\]_sky130_fd_sc_hd__and4_2_B/D
+ VGND VGND VPWR VPWR data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/D sky130_fd_sc_hd__and4_1
Xm_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout161/X m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout614/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_48_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_23_clk_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_845 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_19_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[10\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold667/X hold541/X fanout566/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_38_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A hold1260/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout603/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X
+ m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B fanout394/X fanout238/X
+ m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2/Y VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/A1
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout49/X fanout73/X
+ m_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A_B
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B_A fanout486/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_B1_sky130_fd_sc_hd__or3_2_X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or4_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2/B1
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold324/A m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__and2_2_B/X fanout383/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XANTENNA_fanout113_A fanout115/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__o31ai_2_B1
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2/A1
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/A2
+ sky130_fd_sc_hd__o31ai_4
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold234/A m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__and2_2_B/X fanout396/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.g_buffer\[25\].m_y_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[4\]_sky130_fd_sc_hd__mux2_1_A0 hold457/X m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N/X
+ fanout363/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA_m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__mux2_1_A0_A0 m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout50/X fanout74/X
+ hold1151/A m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_25_1065 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1060/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[2\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1178/X hold1038/X fanout576/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A0 hold46/A m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_S fanout231/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout26_A fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR fanout99/A sky130_fd_sc_hd__and4_2
XFILLER_25_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout155/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B/Y m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_1
XFILLER_36_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold346/A fanout49/X fanout45/X hold1009/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[12\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1031/X m_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout595/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.a0\[2\]_sky130_fd_sc_hd__xnor2_2_Y/A m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X/A2
+ m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B/X
+ sky130_fd_sc_hd__or3b_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold690/A fanout114/X fanout98/X m_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold947/A fanout24/X fanout28/X hold1029/A m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_matrix\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1049/X m_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout562/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold817/X hold1196/A fanout543/X VGND VGND VPWR VPWR hold818/A sky130_fd_sc_hd__mux2_1
XFILLER_79_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__xnor2_2_A m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_37_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__xnor2_1
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_834 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout255/X m_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout373/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold930/X m_blake2.m_hash256.m_matrix\[6\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout588/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_48_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X fanout270/X m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/X
+ m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X/B1 m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X/X sky130_fd_sc_hd__o2bb2a_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__nor2_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout273/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and3_2_A m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B fanout481/X VGND
+ VGND VPWR VPWR fanout420/A sky130_fd_sc_hd__and3_2
Xm_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2_2
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1172/A fanout32/X fanout76/X hold856/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout422/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold693/A fanout26/X m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_2
XANTENNA_m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__o211a_2_X_B1
+ fanout239/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold418 hold418/A VGND VGND VPWR VPWR hold418/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold407 hold407/A VGND VGND VPWR VPWR hold407/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[31\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xhold429 hold429/A VGND VGND VPWR VPWR hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__and3_2_C_B fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__a31o_2_B1 m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ hold1254/A m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__and2_2_A/B
+ m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1 VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_65_1390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_1254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold1129 hold1129/A VGND VGND VPWR VPWR hold1129/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1118 hold1118/A VGND VGND VPWR VPWR hold1118/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold1073/A fanout109/X fanout144/X hold744/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xhold1107 hold1107/A VGND VGND VPWR VPWR hold1107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_61_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[30\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
XFILLER_39_878 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout153/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xtt_um_essen_628 VGND VGND VPWR VPWR tt_um_essen_628/HI uio_out[6] sky130_fd_sc_hd__conb_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout160/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold363/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_61_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_723 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__nor2_2_Y
+ m_io.cmd\[5\]_sky130_fd_sc_hd__and2b_2_B/X m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X
+ VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__nor2_2
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout230_A fanout232/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout328_A fanout330/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__or2_2_B fanout498/X hold23/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_33_1356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_X fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold930 hold930/A VGND VGND VPWR VPWR hold930/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold963 hold963/A VGND VGND VPWR VPWR hold963/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 hold952/A VGND VGND VPWR VPWR hold952/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold941 hold941/A VGND VGND VPWR VPWR hold941/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout199/X m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[172\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout191/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_73_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold974 hold974/A VGND VGND VPWR VPWR hold974/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 hold985/A VGND VGND VPWR VPWR hold985/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold996 hold996/A VGND VGND VPWR VPWR hold996/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout485_X fanout485/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[163\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_1327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold181/X fanout337/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout415/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__xnor2_2_B hold1107/A hold791/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[22\].m_c_buf m_blake2.m_hash256.g_buffer\[22\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[22\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_1250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_1201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[44\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout422/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout146/X
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1 m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/C m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_9_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout196/X m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout189/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y
+ fanout467/X fanout476/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1/B1 sky130_fd_sc_hd__nor2_1
XFILLER_8_215 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__mux2_1_A0 hold316/A m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout384/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout131/X
+ fanout151/X hold649/A m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__and2_2_B fanout439/X hold150/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_10_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold814/X fanout560/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold889/A fanout128/X fanout93/X hold1206/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_0_660 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout359/X m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__a22o_2_A1/X fanout179/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XFILLER_48_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_c_buf\[29\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_c_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_c_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_c_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout175/A hold834/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[29\].m_c_buf/A
+ sky130_fd_sc_hd__o32a_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A0 hold124/A m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[27\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold576/X m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout234/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold119/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__xnor2_2_A hold1086/A hold789/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold893/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2
+ fanout287/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2
+ m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout530/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__mux2_1_A1_S fanout499/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xhash\[7\]_sky130_fd_sc_hd__and2_2_B fanout442/X hash\[7\]_sky130_fd_sc_hd__and2_2_B/B
+ VGND VGND VPWR VPWR hash\[7\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[13\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1199/X m_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout558/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold215 hold215/A VGND VGND VPWR VPWR hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 hold204/A VGND VGND VPWR VPWR hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__and3_2_A hold220/A fanout464/X fanout392/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xhold226 hold226/A VGND VGND VPWR VPWR hold226/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold259/A VGND VGND VPWR VPWR hold259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 hold248/A VGND VGND VPWR VPWR hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 hold237/A VGND VGND VPWR VPWR hold237/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[10\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold456/A sky130_fd_sc_hd__dfxtp_1
XFILLER_63_1327 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
XFILLER_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_c_buf\[1\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or2_2_X
+ hold675/A fanout101/X VGND VGND VPWR VPWR ANTENNA_2/DIODE sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout307/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout180_A fanout180/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A fanout279/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_697 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout244/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__or2_2_B fanout484/X hold137/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold879/X fanout223/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xdata\[0\]_sky130_fd_sc_hd__mux2_1_A1 hold11/X hold9/X fanout598/X VGND VGND VPWR
+ VPWR data\[0\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold394/X m_blake2.m_hash256.v_q\[15\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout211/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold332/A m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout390/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout612_A fanout615/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout233_X fanout233/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_S fanout412/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold385/X m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout158/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold908/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout400_X fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_12_Left_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__inv_2_A m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__inv_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold782 hold782/A VGND VGND VPWR VPWR hold782/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 hold771/A VGND VGND VPWR VPWR hold771/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold760 hold760/A VGND VGND VPWR VPWR hold760/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold708/A fanout83/X fanout67/X hold522/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[9\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold938/X m_blake2.m_hash256.m_matrix\[9\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout603/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout182/X m_blake2.m_hash256.v_q\[4\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_4
Xm_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__a22o_2_A1/X sky130_fd_sc_hd__a22o_1
XFILLER_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold793 hold793/A VGND VGND VPWR VPWR hold793/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold808/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold761/X m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_57_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_d\[25\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1023/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
XTAP_TAPCELL_ROW_4_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_837 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__a21bo_2_B1_N/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ sky130_fd_sc_hd__a21bo_1
Xm_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold117/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_68_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_64_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_531 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1252/X hold917/X fanout577/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout183/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold679/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y
+ fanout347/X m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__nor2_1
XFILLER_40_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold294/X m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout232/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR fanout249/A sky130_fd_sc_hd__or2_4
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout49/X fanout45/X
+ hold917/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold591/A sky130_fd_sc_hd__dfxtp_1
XFILLER_12_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[25\]_sky130_fd_sc_hd__a22o_2_A1_A2 m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1004/X m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout596/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N/X
+ sky130_fd_sc_hd__a21bo_1
Xm_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold551/A fanout96/X fanout120/X hold840/A m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C fanout458/X fanout459/X
+ fanout462/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_buffer\[23\].m_y_buf m_blake2.m_hash256.g_buffer\[23\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[23\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_910 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1
+ fanout363/X m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1/X
+ m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__a211oi_2_A1/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout426/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
XFILLER_36_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_c_buf\[19\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout254/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold431/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__a32o_2_A1 hold1118/A fanout346/X
+ fanout249/X fanout169/X m_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[1\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a32o_1
XFILLER_17_881 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_851 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__and2_2_B fanout430/X hold87/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_50_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_clk_X clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout83/X fanout43/X
+ hold1082/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1
+ fanout427/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A0 hold33/A m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout520/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[49\]_sky130_fd_sc_hd__and3_2_A_B fanout463/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B_A fanout486/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[1\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold968/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold799/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_70_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_67_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout514 fanout515/X VGND VGND VPWR VPWR fanout514/X sky130_fd_sc_hd__clkbuf_4
Xfanout503 fanout504/X VGND VGND VPWR VPWR fanout503/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/Y m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/C
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/B
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold599/X m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B fanout429/X hold51/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xfanout536 fanout537/X VGND VGND VPWR VPWR fanout536/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_fanout395_A fanout398/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout547 fanout548/X VGND VGND VPWR VPWR fanout547/X sky130_fd_sc_hd__clkbuf_4
Xfanout525 fanout526/X VGND VGND VPWR VPWR fanout525/X sky130_fd_sc_hd__clkbuf_4
Xfanout558 fanout561/X VGND VGND VPWR VPWR fanout558/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout569 fanout570/X VGND VGND VPWR VPWR fanout569/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout183_X fanout183/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_6_1051 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X_B1 m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout350_X fanout350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout19/X m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[27\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XANTENNA_fanout448_X fanout448/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[10\]\[6\]_sky130_fd_sc_hd__mux2_1_A0 hold671/X m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[5\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1248/X m_blake2.m_hash256.m_matrix\[6\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout581/X
+ VGND VGND VPWR VPWR hold1249/A sky130_fd_sc_hd__mux2_1
XFILLER_42_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold369/A fanout34/X fanout74/X hold1115/A m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[3\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold957/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout615_X fanout615/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold610/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_Q hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold705/A fanout138/X fanout95/X hold319/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/Y sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B
+ fanout254/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold79/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[115\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold600/X fanout326/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold964/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X/A1
+ fanout368/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2
+ sky130_fd_sc_hd__nand2_8
XFILLER_11_1292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y
+ fanout446/X m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR hold217/A sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout348/X m_blake2.m_hash256.v_q\[5\]\[19\]_sky130_fd_sc_hd__a22o_2_A1/X fanout178/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_57_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B fanout498/X hold113/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[239\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xhold590 hold590/A VGND VGND VPWR VPWR hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout96_X fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold305/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.g_buffer\[27\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[14\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A fanout454/X fanout456/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/C VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__inv_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A0 hold140/A m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout504/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[8\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1084/A fanout48/X fanout68/X hold780/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[3\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1005/X hold954/X fanout600/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout153/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_781 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__o21bai_2_A1/Y m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1/X
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__or4_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold309/A sky130_fd_sc_hd__dfxtp_1
XFILLER_36_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X
+ hold976/A fanout143/X fanout95/X m_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_19_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold956/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_832 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_865 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A/B m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_fanout310_A fanout314/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout408_A fanout408/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__a22o_2_A1 hold713/X fanout339/X
+ m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__a22o_2_A1/B1 fanout535/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout357/X m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X fanout257/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold392/X m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B
+ fanout329/X m_blake2.m_hash256.h_flat\[140\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[8\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.v_q\[8\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1091/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[1\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1242/X hold1252/A fanout575/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout322 fanout323/X VGND VGND VPWR VPWR fanout322/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout621/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout398_X fanout398/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout311 fanout312/X VGND VGND VPWR VPWR fanout311/X sky130_fd_sc_hd__clkbuf_4
Xfanout300 fanout301/X VGND VGND VPWR VPWR fanout300/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload21/A m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_1113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[22\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
Xfanout344 fanout345/X VGND VGND VPWR VPWR fanout344/X sky130_fd_sc_hd__dlymetal6s2s_1
Xfanout333 fanout334/X VGND VGND VPWR VPWR fanout333/X sky130_fd_sc_hd__clkbuf_4
Xfanout355 fanout361/X VGND VGND VPWR VPWR fanout355/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1/B1 m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_6_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__o22a_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout366 fanout371/X VGND VGND VPWR VPWR fanout366/X sky130_fd_sc_hd__buf_2
XFILLER_74_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout399 fanout399/A VGND VGND VPWR VPWR fanout399/X sky130_fd_sc_hd__buf_4
Xfanout377 fanout399/X VGND VGND VPWR VPWR fanout377/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
Xfanout388 fanout391/X VGND VGND VPWR VPWR fanout388/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/A2
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1256/X m_blake2.m_hash256.m_matrix\[11\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout591/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold696/A fanout126/X fanout114/X hold1222/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.g_d\[31\]_sky130_fd_sc_hd__o21a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[8\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1136/X hold1123/X fanout551/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_35_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_858 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[30\]_sky130_fd_sc_hd__a22o_2_X_A1 fanout355/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_1376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold1015/A fanout57/X fanout69/X hold566/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[8\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[27\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.res_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/A fanout260/X
+ m_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__a221o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_A
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X hold277/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[5\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.fsm_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
XFILLER_19_965 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.h_flat\[242\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold224/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_29_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X
+ m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[121\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold225/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold741/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout169/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_1243 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold212/X fanout316/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X_sky130_fd_sc_hd__a21o_2_A2
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A2
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout182/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__xnor2_2_A hold419/A hold1218/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__a22o_2_A1 hold428/A fanout290/X
+ fanout278/X hold524/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ fanout450/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/B
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__and2_2_B fanout433/X hold615/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/A
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/B
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/A
+ sky130_fd_sc_hd__and3_1
XFILLER_60_1105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a2111o_2_A2
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C/X
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1/X
+ m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a2111o_2_A2/X
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_9_1433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_27_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_902 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout260_A fanout265/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout358_A fanout361/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_1045 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1034 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__xnor2_2_B hold1110/A hold452/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_75_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout146_X fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_S fanout412/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_684 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__xnor2_2_A hold358/A hold819/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold867/X hold1201/A fanout565/X VGND VGND VPWR VPWR hold868/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__or2_2_B fanout498/X hold17/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout419/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold319/X fanout606/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_3_6_0_clk_X clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout130 fanout131/A VGND VGND VPWR VPWR fanout130/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout163 fanout168/A VGND VGND VPWR VPWR fanout163/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold167/A sky130_fd_sc_hd__dfxtp_1
Xfanout152 fanout152/A VGND VGND VPWR VPWR fanout152/X sky130_fd_sc_hd__buf_2
XFILLER_43_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout141 fanout143/X VGND VGND VPWR VPWR fanout141/X sky130_fd_sc_hd__buf_2
Xfanout174 fanout174/A VGND VGND VPWR VPWR fanout174/X sky130_fd_sc_hd__clkbuf_8
Xfanout196 fanout197/X VGND VGND VPWR VPWR fanout196/X sky130_fd_sc_hd__clkbuf_4
Xfanout185 fanout186/A VGND VGND VPWR VPWR fanout185/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B/X
+ sky130_fd_sc_hd__and3b_1
XFILLER_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__and2_2_B_A fanout442/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[156\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold26/X fanout329/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout587/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold168/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[2\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold152/X fanout325/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B fanout434/X hold136/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[52\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_11_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__xnor2_2_A hold703/A hold858/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__and2_2_B fanout433/X hold632/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1079/A fanout84/X fanout120/X hold549/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout182/X m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_4
XPHY_EDGE_ROW_0_Left_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout101/X hold1233/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o32a_2
Xm_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X m_io.m_config.ll_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold204/A sky130_fd_sc_hd__dfxtp_1
XFILLER_66_857 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__a211o_2_A1 hold789/A fanout293/X
+ m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__a22o_2_A1/X fanout390/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[7\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A0 hold36/A m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout512/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[12\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1227/X hold1155/X fanout558/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1220/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_743 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_765 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__xnor2_2_A hold396/A hold940/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_hash\[2\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2_A1 fanout401/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_hash\[2\]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2_B2 fanout285/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[249\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout195/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__and3_2_B m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__xnor2_2_B hold1046/A hold411/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold961/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1_C1 m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout106_A fanout107/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_8_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_1336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold863/A fanout87/X fanout135/X hold563/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold195/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout475_A fanout476/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__xnor2_2_A hold393/A hold907/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XFILLER_25_1077 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0 hold356/A hash\[7\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout391/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold46/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_38_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout430_X fanout430/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout246/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_43_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[8\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold983/X hold790/X fanout600/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_37_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.g_buffer\[31\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1 hold510/A fanout278/X
+ m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__a22o_2_A1/X fanout367/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout80/X
+ fanout64/X m_blake2.m_hash256.m_matrix\[11\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[19\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A0_S fanout520/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A0 hold261/A m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_S fanout213/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[41\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N
+ m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold643/X fanout165/X m_io.m_config.ll_q\[23\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X
+ hold624/A fanout87/X fanout119/X hold1158/A m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a221o_1
Xhold408 hold408/A VGND VGND VPWR VPWR hold408/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 hold419/A VGND VGND VPWR VPWR hold419/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_61_1222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_61_1233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X hold255/X
+ fanout163/X m_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__or2_2_A/X fanout616/X VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout198/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1108 hold1108/A VGND VGND VPWR VPWR hold1108/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1119 hold1119/A VGND VGND VPWR VPWR hold1119/X sky130_fd_sc_hd__dlygate4sd3_1
Xtt_um_essen_629 VGND VGND VPWR VPWR tt_um_essen_629/HI uio_out[5] sky130_fd_sc_hd__conb_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[26\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
XFILLER_80_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1026 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__xnor2_2_A hold1037/A hold792/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_22_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_33_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_779 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold142/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
XANTENNA_fanout223_A fanout224/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold931 hold931/A VGND VGND VPWR VPWR hold931/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold920 hold920/A VGND VGND VPWR VPWR hold920/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 hold964/A VGND VGND VPWR VPWR hold964/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 hold942/A VGND VGND VPWR VPWR hold942/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X
+ hold764/A fanout146/X fanout122/X hold1164/A m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/A2
+ sky130_fd_sc_hd__a221o_1
Xhold953 hold953/A VGND VGND VPWR VPWR hold953/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold986 hold986/A VGND VGND VPWR VPWR hold986/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 hold997/A VGND VGND VPWR VPWR hold997/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold975 hold975/A VGND VGND VPWR VPWR hold975/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__or3_2_B_A fanout407/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[4\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1115/X hold1222/A fanout580/X VGND VGND VPWR VPWR hold1116/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout478_X fanout478/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold257/X fanout166/X m_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_40_1317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold55/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_45_849 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_77_1262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ hold652/X m_io.m_config.cfg_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o21a_1
XFILLER_71_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_724 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold286/A sky130_fd_sc_hd__dfxtp_1
XFILLER_44_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[26\].m_c_buf m_blake2.m_hash256.g_buffer\[26\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[26\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_22_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_B1 fanout401/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__xor2_2_A hold463/A hold367/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_10_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[63\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_39_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_37_clk_A clkload5/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__or2_2_B fanout485/X hold32/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[145\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold264/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[12\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold348/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[10\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold365/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2_A1
+ hash\[4\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_952 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold353/A fanout126/X fanout86/X hold1094/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[189\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold124/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[12\]\[5\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold831/X fanout227/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_36_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ hold505/X fanout305/X m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
XANTENNA_clkload1_A clkload1/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout85/X fanout113/X
+ hold1080/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold652/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[2\]_sky130_fd_sc_hd__a211o_2_X_A1 m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold1019/X m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold876/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[2\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold873/X hold811/X fanout574/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold963/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and2_2_B fanout430/X hold164/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xhold216 hold216/A VGND VGND VPWR VPWR hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 hold205/A VGND VGND VPWR VPWR hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A VGND VGND VPWR VPWR hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[12\]\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/B fanout227/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1112/A fanout88/X fanout149/X hold654/A m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xhold249 hold249/A VGND VGND VPWR VPWR hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 hold227/A VGND VGND VPWR VPWR hold227/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_67_1453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_63_1339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[2\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold780/X fanout571/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A hold3/X m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_61_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[15\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold752/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_1172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/A1
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/A3
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nand2_1
XFILLER_6_1244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_1003 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[12\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold955/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout183/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.m_matrix\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold863/X hold839/X fanout601/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout173_A fanout173/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B_A fanout487/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold338/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout340_A fanout341/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_A
+ fanout269/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/A1 hold897/X fanout577/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout438_A fanout442/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__or2_2_B fanout491/X hold33/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold332/X fanout412/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a22o_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/A sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_20_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0 hold459/X m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X/B2
+ fanout556/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ fanout237/X m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/X m_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X
+ fanout270/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__mux2_1_A0_S fanout520/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[10\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout593/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout182/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold460/A sky130_fd_sc_hd__dfxtp_1
Xhold772 hold772/A VGND VGND VPWR VPWR hold772/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold750 hold750/A VGND VGND VPWR VPWR hold750/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold761 hold761/A VGND VGND VPWR VPWR hold761/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_io.m_config.ll_q\[63\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold794 hold794/A VGND VGND VPWR VPWR hold794/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout86_A fanout87/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold783 hold783/A VGND VGND VPWR VPWR hold783/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_77_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_58_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1027/X hold1208/A fanout543/X VGND VGND VPWR VPWR hold1028/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_45_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout283/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_849 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_808 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_819 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold275/X m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout210/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_882 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[4\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold370/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_64_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_A
+ fanout473/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold322/A m_blake2.m_hash256.h_flat\[202\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout370/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_885 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or3b_2_B/C_N
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X
+ fanout269/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold771/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold569/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_1345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_63_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[27\].m_y_buf m_blake2.m_hash256.g_buffer\[27\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[27\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[19\]_sky130_fd_sc_hd__o22a_2_X_A2 fanout175/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_1130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold125/A sky130_fd_sc_hd__dfxtp_1
XFILLER_56_1110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout193/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[224\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold33/X fanout327/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[216\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
XTAP_TAPCELL_ROW_14_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout120/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold416/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_3_7_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload5/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__a22o_2_A1_A1 m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkload21/A m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold792/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X
+ hold725/A fanout139/X fanout107/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y
+ fanout469/X m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_70_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout515 fanout516/X VGND VGND VPWR VPWR fanout515/X sky130_fd_sc_hd__clkbuf_4
Xfanout504 fanout509/X VGND VGND VPWR VPWR fanout504/X sky130_fd_sc_hd__buf_2
Xfanout537 fanout538/X VGND VGND VPWR VPWR fanout537/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_738 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y
+ fanout184/X m_blake2.m_hash256.v_q\[4\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1/X m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y/A sky130_fd_sc_hd__o21ai_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_A_N
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout548 fanout550/X VGND VGND VPWR VPWR fanout548/X sky130_fd_sc_hd__clkbuf_4
Xfanout526 fanout538/X VGND VGND VPWR VPWR fanout526/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout559 fanout560/X VGND VGND VPWR VPWR fanout559/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout290_A fanout291/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_X fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold716/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout450/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold709/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_646 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout231/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[5\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold931/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_14_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__xnor2_2_A hold655/A hold1220/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_39_1352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__a21o_2_X/A2
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/B sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_25_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold1050/A fanout56/X fanout68/X hold1146/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3
+ fanout451/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3/X
+ sky130_fd_sc_hd__o31a_1
Xm_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A0 hold211/A m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X/B sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_12_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout608_X fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__mux2_1_A0 hold157/A m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout518/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1009 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold580 hold580/A VGND VGND VPWR VPWR hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[7\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold758/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X_B2_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[13\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1169/A hold1029/X fanout559/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold591 hold591/A VGND VGND VPWR VPWR hold591/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_C1
+ fanout268/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__xor2_2_B hold448/A hold384/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1 m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/C m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_79_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_io.cmd\[2\]_sky130_fd_sc_hd__o21ai_2_A1 block_last_sky130_fd_sc_hd__a32o_2_B2/A1
+ block_last_sky130_fd_sc_hd__a32o_2_B2/A2 block_last_sky130_fd_sc_hd__a32o_2_B2/A3
+ VGND VGND VPWR VPWR fanout308/A sky130_fd_sc_hd__o21ai_2
XTAP_TAPCELL_ROW_66_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_402 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[10\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold994/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold395/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_947 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X
+ hold976/A fanout27/X m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a2111o_1
Xm_blake2.m_hash256.m_matrix\[9\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold880/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[14\]_sky130_fd_sc_hd__a2bb2o_2_A1_N hold547/A fanout380/X
+ fanout264/X hold1008/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1/B1
+ sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_2
XANTENNA_m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__and3_2_C_A fanout448/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold140/X fanout312/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[34\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold608/X m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1 hold932/A fanout351/X
+ fanout263/X m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[38\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N
+ fanout418/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1/X
+ VGND VGND VPWR VPWR fanout299/A sky130_fd_sc_hd__o21ba_2
Xm_blake2.m_hash256.m_matrix\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[5\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1080/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_B1
+ fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1125/X m_blake2.m_hash256.m_matrix\[12\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout565/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout200/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout258/X m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ fanout381/X fanout180/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ hold371/A fanout306/X m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__mux2_1_A0 hold123/A m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X m_io.m_config.ll_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold573/A sky130_fd_sc_hd__dfxtp_1
XFILLER_52_903 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_S fanout418/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A0 hold188/A m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_958 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout136_A fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A0 hold38/A m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_899 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout303_A fanout303/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout323 fanout342/A VGND VGND VPWR VPWR fanout323/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_2
Xfanout301 fanout303/A VGND VGND VPWR VPWR fanout301/X sky130_fd_sc_hd__clkbuf_4
Xfanout312 fanout314/X VGND VGND VPWR VPWR fanout312/X sky130_fd_sc_hd__buf_2
Xfanout345 fanout346/X VGND VGND VPWR VPWR fanout345/X sky130_fd_sc_hd__buf_2
Xfanout356 fanout361/X VGND VGND VPWR VPWR fanout356/X sky130_fd_sc_hd__buf_2
Xfanout334 fanout335/X VGND VGND VPWR VPWR fanout334/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout367 fanout371/X VGND VGND VPWR VPWR fanout367/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold98/A sky130_fd_sc_hd__dfxtp_1
Xfanout389 fanout391/X VGND VGND VPWR VPWR fanout389/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1 hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout378 fanout379/X VGND VGND VPWR VPWR fanout378/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_matrix\[7\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold520/X hold821/A fanout602/X VGND VGND VPWR VPWR hold521/A sky130_fd_sc_hd__mux2_1
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout49_A fanout51/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_A1
+ fanout288/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_B2
+ fanout283/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1095 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_2_0_clk_X clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_Y
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_1418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_55_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__o211a_2_A1 m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__o211a_2_A1/X sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B fanout497/X hold195/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__mux2_1_A1_S fanout223/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold462/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__nand2_2_Y
+ m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_io.m_config.ll_q\[41\]_sky130_fd_sc_hd__and3_2_A_B fanout463/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[18\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout188/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2/A1
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_2
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand3_2_C/B
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout232/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_741 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A0 hold177/A m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_2
XFILLER_18_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_1293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_40_clk clkload5/A VGND VGND VPWR VPWR clkbuf_leaf_40_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_41_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_69_822 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__a21oi_2_B1 m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_37_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_2
XFILLER_25_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout253_A fanout254/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_917 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout139_X fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clkload4/A VGND VGND VPWR VPWR clkload30/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__nor2_2_B fanout495/X hold184/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout420_A fanout420/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR fanout147/A sky130_fd_sc_hd__and4_2
Xm_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1151/X fanout581/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__mux2_1_A0 hold1150/X m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__xor2_2_A hold580/A hold808/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1149/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A2
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1/Y
+ sky130_fd_sc_hd__o211ai_1
Xm_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_50_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout131 fanout131/A VGND VGND VPWR VPWR fanout131/X sky130_fd_sc_hd__clkbuf_2
Xfanout120 fanout123/X VGND VGND VPWR VPWR fanout120/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__xnor2_2_A hold440/A hold1024/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xfanout164 fanout168/X VGND VGND VPWR VPWR fanout164/X sky130_fd_sc_hd__buf_2
Xfanout142 fanout143/X VGND VGND VPWR VPWR fanout142/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__a31o_2_B1 m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[28\]_sky130_fd_sc_hd__and2_2_A/B
+ m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.block_idx_plus_one_q\[30\]_sky130_fd_sc_hd__a31o_2_B1/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_1 fanout454/X fanout456/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C/X m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_1/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout153 fanout154/X VGND VGND VPWR VPWR fanout153/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold984/A fanout84/X fanout113/X hold853/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__a2bb2o_2_A1_N hold391/A fanout382/X
+ fanout264/X m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__a2bb2o_2_A1_N/B2
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/B1 sky130_fd_sc_hd__a2bb2o_1
Xfanout197 fanout200/A VGND VGND VPWR VPWR fanout197/X sky130_fd_sc_hd__buf_2
Xfanout186 fanout186/A VGND VGND VPWR VPWR fanout186/X sky130_fd_sc_hd__clkbuf_4
XFILLER_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_S fanout156/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout175 fanout175/A VGND VGND VPWR VPWR fanout175/X sky130_fd_sc_hd__buf_4
XFILLER_19_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_S fanout160/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout288/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_733 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__xnor2_2_B hold1137/A hold466/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_70_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout343/X m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ fanout177/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a211o_1
XFILLER_54_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_22_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkload16/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__xnor2_2_A hold964/A hold532/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_667 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__xor2_2_A hold305/A hold707/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XFILLER_13_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_803 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold86/A sky130_fd_sc_hd__dfxtp_1
XFILLER_65_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[1\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold772/X hold947/X fanout574/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold36/X fanout320/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X
+ fanout239/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1/Y
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_4_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_1 hold256/A m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout397/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout245/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_55_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
Xclkbuf_leaf_13_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_13_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_io.hash_v_o_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X hash_v_sky130_fd_sc_hd__a211o_2_X/X
+ VGND VGND VPWR VPWR uio_out_sky130_fd_sc_hd__buf_2_X_1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_31_1274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1266/A fanout128/X fanout144/X m_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_66_1315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout88/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__xnor2_2_A hold232/A hold1210/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A_A fanout472/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__or3b_2_A/B fanout481/X VGND
+ VGND VPWR VPWR fanout412/A sky130_fd_sc_hd__or3b_4
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_S fanout233/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[14\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold339/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout370_A fanout371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A0 hold1061/A m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout520/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_80_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout256_X fanout256/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__xnor2_2_A hold956/A hold538/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_A1 fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__mux2_1_A1_S fanout489/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_1065 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[204\]_sky130_fd_sc_hd__or2_2_B_A fanout499/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold615/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1051/X fanout545/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold975/A fanout132/X fanout136/X m_blake2.m_hash256.m_matrix\[2\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_37_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[8\]\[25\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ fanout355/X fanout253/X VGND VGND VPWR VPWR fanout175/A sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold253/A sky130_fd_sc_hd__dfxtp_1
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout194/X m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[14\]\[30\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout176/X fanout272/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1/X m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/A3
+ m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2/X
+ sky130_fd_sc_hd__a31o_2
Xm_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[6\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XFILLER_48_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_817 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold261/X fanout325/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1005/A fanout56/X fanout46/X hold873/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1020/A fanout112/X fanout137/X hold969/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__nand2_2_B fanout434/X hold154/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[84\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__a22o_2_A1 hold501/A fanout294/X
+ fanout286/X hold681/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ fanout344/X m_blake2.m_hash256.h_flat\[234\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X fanout255/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__mux2_1_A0 hold439/A m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout367/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__o311a_2_A1 m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/A
+ hold1217/A m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/Y fanout308/A
+ fanout611/X VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__o311a_2_A1/X
+ sky130_fd_sc_hd__o311a_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/B2
+ m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout274/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o22a_1
Xm_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[3\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
XFILLER_16_766 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_714 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A1_S fanout411/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__and3b_2_X
+ fanout475/X fanout469/X fanout466/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ sky130_fd_sc_hd__and3b_4
XFILLER_54_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold409 hold409/A VGND VGND VPWR VPWR hold409/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[24\]_sky130_fd_sc_hd__or2_2_A hold986/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[24\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_48_1001 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[13\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold748/X m_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout563/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__or2_2_B fanout483/X hold274/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A0 hold192/A m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout512/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold1110/X m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout233/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ hold1255/X m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout426/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[55\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1164/X
+ fanout583/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__a22o_2_A1 hold336/A fanout190/X
+ fanout198/X hold670/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold656/X fanout606/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1 m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR fanout258/A sky130_fd_sc_hd__or2_4
Xhold1109 hold1109/A VGND VGND VPWR VPWR hold1109/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[3\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold693/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_2_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkload6/A sky130_fd_sc_hd__clkbuf_8
XFILLER_66_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__or2_2_A hold1062/A fanout367/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_0_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__a22o_2_A1 hold756/A fanout188/X
+ fanout196/X hold875/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[10\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ hold913/X VGND VGND VPWR VPWR hold912/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_77_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold921 hold921/A VGND VGND VPWR VPWR hold921/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold910 hold910/A VGND VGND VPWR VPWR hold910/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 hold932/A VGND VGND VPWR VPWR hold932/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold954 hold954/A VGND VGND VPWR VPWR hold954/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold943 hold943/A VGND VGND VPWR VPWR hold943/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout160/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold987 hold987/A VGND VGND VPWR VPWR hold987/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold965 hold965/A VGND VGND VPWR VPWR hold965/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold976 hold976/A VGND VGND VPWR VPWR hold976/X sky130_fd_sc_hd__dlygate4sd3_1
Xdata\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X data\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold179/A sky130_fd_sc_hd__dfxtp_1
Xhold998 hold998/A VGND VGND VPWR VPWR hold998/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_27_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold389/X m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[12\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold445/A sky130_fd_sc_hd__dfxtp_1
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata\[5\]_sky130_fd_sc_hd__mux2_1_A1 data\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold1047/X
+ fanout550/X VGND VGND VPWR VPWR data\[5\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_32_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1021/A sky130_fd_sc_hd__dfxtp_1
XFILLER_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_1214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold900/A fanout84/X fanout116/X hold1250/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__xor2_2_B/A fanout219/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout82/X
+ fanout42/X hold1072/A m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B/A
+ fanout407/X VGND VGND VPWR VPWR fanout288/A sky130_fd_sc_hd__nor2_8
Xm_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold1098/A fanout275/X fanout176/X m_blake2.m_hash256.v_q\[14\]\[13\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout272/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_60_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1039/X m_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout578/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_23_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_10_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold696/X m_blake2.m_hash256.m_matrix\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout581/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_39_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_5_979 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[2\]_sky130_fd_sc_hd__mux2_1_A1_S fanout205/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold915/X fanout208/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o211a_2_A2_C1
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold464/X m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout258/X m_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout382/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__a22o_2_A1/B1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_36_839 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__xnor2_2_B hold281/A hold524/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__xnor2_2_B/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold572/A sky130_fd_sc_hd__dfxtp_1
XFILLER_62_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_Q hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21a_2_A1
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__o21a_1
XANTENNA_block_first_sky130_fd_sc_hd__a22o_2_B2_A1 fanout485/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__and3_2_A hold257/A fanout464/X fanout392/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XFILLER_56_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold398/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1063/X
+ fanout565/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0 hold318/X m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout420/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_31_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_28_Left_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[18\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold206 hold206/A VGND VGND VPWR VPWR hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold217/A VGND VGND VPWR VPWR hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold228 hold228/A VGND VGND VPWR VPWR hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 hold239/A VGND VGND VPWR VPWR hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__and2_2
XFILLER_67_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1113/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout295/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_37_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold507/X m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1075 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold1039/A fanout83/X fanout74/X m_blake2.m_hash256.m_matrix\[4\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__a32o_2_A1_B1 fanout170/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold753/X m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR
+ VPWR hold134/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_46_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[13\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1053/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_79_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout500_A fanout500/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A1
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__or3_2_C/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/A
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1060/A fanout134/X fanout94/X hold1090/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[0\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[0\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold453/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[6\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold722/X hold992/A fanout573/X VGND VGND VPWR VPWR hold723/A sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold303/X fanout165/X m_io.m_config.ll_q\[21\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_2_916 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[48\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[47\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_55_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y
+ fanout220/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[26\]_sky130_fd_sc_hd__a211o_2_X hold941/A fanout174/X
+ m_blake2.m_hash256.g_c_buf\[26\]_sky130_fd_sc_hd__a211o_2_X/B1 m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__a32o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[26\].m_c_buf/A sky130_fd_sc_hd__a211o_1
Xhold773 hold773/A VGND VGND VPWR VPWR hold773/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold762 hold762/A VGND VGND VPWR VPWR hold762/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 hold751/A VGND VGND VPWR VPWR hold751/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold740 hold740/A VGND VGND VPWR VPWR hold740/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 hold795/A VGND VGND VPWR VPWR hold795/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__a21bo_2_B1_N/X m_blake2.m_hash256.m_g.m_add_1.x2_i\[19\]_sky130_fd_sc_hd__nand3b_2_A_N/Y
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/C
+ sky130_fd_sc_hd__a21o_1
Xhold784 hold784/A VGND VGND VPWR VPWR hold784/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_39_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_S fanout153/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[15\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold886/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__or2_2_A hold226/A fanout380/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_4_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold904/X m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout155/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_68_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold873/A sky130_fd_sc_hd__dfxtp_1
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_64_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout34_X fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1/B1
+ sky130_fd_sc_hd__inv_2
XFILLER_38_1022 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A1 m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_64_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold322/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_71_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1
+ m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1/Y
+ VGND VGND VPWR VPWR fanout160/A sky130_fd_sc_hd__nor2_2
XFILLER_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_B
+ fanout477/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B
+ fanout426/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1/X m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_73_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold710/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[4\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1108/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout347/X m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__a22o_2_A1/X fanout177/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout195/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[8\]\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold726/X fanout224/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_1357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_4
XFILLER_64_956 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A0 hold88/A m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout529/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold511/X fanout167/X m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__or2_2_A/X fanout618/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_63_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_842 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__a21oi_2_B1 m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[2\]_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[6\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold551/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__o211a_2_A1 m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__o211a_2_A1/X sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold299/A m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__and2_2_B/X fanout376/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__inv_2_Y_A
+ fanout478/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout505 fanout509/X VGND VGND VPWR VPWR fanout505/X sky130_fd_sc_hd__clkbuf_4
Xfanout538 fanout539/X VGND VGND VPWR VPWR fanout538/X sky130_fd_sc_hd__clkbuf_4
Xfanout516 fanout539/X VGND VGND VPWR VPWR fanout516/X sky130_fd_sc_hd__clkbuf_2
Xfanout527 fanout529/X VGND VGND VPWR VPWR fanout527/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_63_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ hold565/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xfanout549 fanout550/X VGND VGND VPWR VPWR fanout549/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1_A1 m_blake2.m_hash256.m_g.d_q\[20\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout283_A fanout283/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1_1/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3/B1
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold1220/X fanout222/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[2\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1096/X hold1153/A fanout556/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout280/X m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout287/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_1_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[21\]_sky130_fd_sc_hd__a221o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[221\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold206/A sky130_fd_sc_hd__dfxtp_1
XFILLER_54_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout169_X fanout169/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X fanout610/X
+ m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X/B VGND VGND
+ VPWR VPWR m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_36_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold931/A fanout39/X fanout47/X hold705/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.h_flat\[100\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold99/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_12_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold211/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_41_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[109\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold157/X fanout325/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__nor2_2_B fanout499/X hold139/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold784/X fanout564/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_57_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold581 hold581/A VGND VGND VPWR VPWR hold581/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold570 hold570/A VGND VGND VPWR VPWR hold570/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1 hold381/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/A2 fanout426/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_57_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold592 hold592/A VGND VGND VPWR VPWR hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_768 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_53_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y
+ m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold853/X hold1070/A fanout568/X VGND VGND VPWR VPWR hold854/A sky130_fd_sc_hd__mux2_1
XFILLER_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1270 hold1270/A VGND VGND VPWR VPWR hold1270/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_input11_A uio_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_66_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold725/X hold705/A fanout605/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold1227/A fanout93/X m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout105/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A1_S fanout411/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_831 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__xnor2_2_A hold316/A hold457/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1/Y m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
XFILLER_9_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1085 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold683/X hold802/A fanout578/X VGND VGND VPWR VPWR hold684/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold886/A fanout61/X fanout37/X hold736/A m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/A m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_B2 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/X fanout609/X input10/X VGND VGND VPWR VPWR m_io.m_config.data_i\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_A1_N
+ fanout188/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold176/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_B1
+ fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold49/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold762/A fanout132/X fanout92/X hold1152/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold853/A fanout37/X fanout45/X hold1259/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_937 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[135\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold188/X fanout333/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__a22o_2_A1 hold677/A fanout292/X
+ fanout286/X hold498/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_71_1428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold38/X fanout314/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_1283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout129_A fanout131/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X m_blake2.m_hash256.g_buffer\[4\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[4\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout498_A fanout499/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout176/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout302 fanout303/X VGND VGND VPWR VPWR fanout302/X sky130_fd_sc_hd__buf_4
Xfanout313 fanout314/X VGND VGND VPWR VPWR fanout313/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_input3_A ui_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout346 fanout361/A VGND VGND VPWR VPWR fanout346/X sky130_fd_sc_hd__clkbuf_4
Xfanout357 fanout361/X VGND VGND VPWR VPWR fanout357/X sky130_fd_sc_hd__buf_2
Xfanout335 fanout342/X VGND VGND VPWR VPWR fanout335/X sky130_fd_sc_hd__buf_4
XTAP_TAPCELL_ROW_6_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout324 fanout325/X VGND VGND VPWR VPWR fanout324/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout368 fanout369/X VGND VGND VPWR VPWR fanout368/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout286_X fanout286/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout379 fanout385/X VGND VGND VPWR VPWR fanout379/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__mux2_1_A0 hold139/A m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout531/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or3_2_C_A
+ fanout346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold307/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_76_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold700/X hold778/A fanout553/X VGND VGND VPWR VPWR hold701/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B
+ m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout530/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X_A2
+ fanout139/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__xnor2_2_A hold332/A hold1191/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_hash\[5\]_sky130_fd_sc_hd__mux2_1_A1_X hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout183/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/X
+ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_46_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1047 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout237/X m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
XFILLER_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[17\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1
+ m_blake2.m_hash256.m_g.d_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or2_2_A fanout461/A fanout462/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/C sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_59_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold958/A fanout86/X fanout110/X m_blake2.m_hash256.m_matrix\[7\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_59_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__a211o_2_A1 hold791/A fanout288/X
+ m_blake2.m_hash256.v_q\[1\]\[5\]_sky130_fd_sc_hd__a22o_2_A1/X fanout379/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout353/X m_blake2.m_hash256.v_q\[5\]\[14\]_sky130_fd_sc_hd__a22o_2_A1/X fanout180/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout292/X m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ fanout356/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2
+ fanout256/X m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.h_flat\[251\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ fanout375/X fanout178/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold137/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ fanout499/X m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_3_6_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload4/A sky130_fd_sc_hd__clkbuf_8
XFILLER_24_1463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[74\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold177/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[66\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_29_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XFILLER_33_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_B2
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__and2_2_B fanout430/X hold474/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__xnor2_2_A hold294/A hold1234/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XFILLER_14_694 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1117/X hold1074/X fanout583/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[67\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[3\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[75\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_31_1401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1 hold942/A fanout348/X
+ fanout260/X m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__or2_2_A hold240/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A0 hold651/A m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout533/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A
+ m_blake2.m_hash256.g_buffer\[10\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold879/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout196/X m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout188/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_3_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__o21ai_2_A1/A2 m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A0 hold122/A m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout36/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__and4_2_C/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_36_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_4
Xm_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold234/X m_blake2.m_hash256.v_q\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout232/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout214/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__xnor2_2_B hold1062/A hold611/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold490/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_2
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR fanout143/A sky130_fd_sc_hd__and4_1
XANTENNA_fanout413_A fanout414/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_664 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold377/X m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_41_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout201_X fanout201/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__xnor2_2_A hold546/A hold831/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[15\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold948/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X/A
+ sky130_fd_sc_hd__and3_1
Xfanout110 fanout111/A VGND VGND VPWR VPWR fanout110/X sky130_fd_sc_hd__clkbuf_4
Xfanout121 fanout123/X VGND VGND VPWR VPWR fanout121/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_S fanout234/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout165 fanout166/X VGND VGND VPWR VPWR fanout165/X sky130_fd_sc_hd__buf_2
Xfanout143 fanout143/A VGND VGND VPWR VPWR fanout143/X sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_50_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout154 fanout156/A VGND VGND VPWR VPWR fanout154/X sky130_fd_sc_hd__clkbuf_4
Xfanout132 fanout135/A VGND VGND VPWR VPWR fanout132/X sky130_fd_sc_hd__clkbuf_4
Xfanout176 fanout176/A VGND VGND VPWR VPWR fanout176/X sky130_fd_sc_hd__buf_4
Xfanout187 fanout189/X VGND VGND VPWR VPWR fanout187/X sky130_fd_sc_hd__clkbuf_4
Xfanout198 fanout200/A VGND VGND VPWR VPWR fanout198/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold415/A fanout112/X fanout140/X m_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_75_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[11\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold503/X m_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout574/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout61_A fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__and3_2_C fanout447/X fanout480/X
+ hold173/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2/X
+ sky130_fd_sc_hd__o21ba_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_48_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_981 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_B1 fanout16/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_A_sky130_fd_sc_hd__and3_2_X
+ fanout467/X fanout469/X fanout474/X VGND VGND VPWR VPWR fanout445/A sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A0 hold115/A m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/A
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ hold291/A fanout306/X m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y/B sky130_fd_sc_hd__a21oi_1
XFILLER_61_1405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_blake2.m_hash256.fsm_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1075/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1160/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1011/A fanout28/X fanout36/X hold415/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_C1
+ fanout346/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload23/A m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[5\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_77_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_B1
+ fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X/A2 m_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[3\].m_c_buf/A sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold811/A fanout136/X fanout144/X m_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold378/A fanout24/X fanout48/X m_blake2.m_hash256.m_matrix\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_18_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout523/X m_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XFILLER_18_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ hold516/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 fanout240/A hold196/A
+ m_blake2.m_hash256.v_q\[12\]\[30\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1_A1 m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1
+ fanout400/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2
+ fanout266/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold747/A fanout33/X fanout69/X m_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[7\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__nor2_2_A_B fanout476/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[69\]_sky130_fd_sc_hd__or2_2_B_A fanout494/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout196_A fanout197/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold543/A fanout44/X fanout72/X hold1108/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X_X m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[168\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold1061/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[160\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1423 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__and3_2_C fanout448/X fanout479/X
+ hold149/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XFILLER_52_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold898/X hold1195/A fanout559/X VGND VGND VPWR VPWR hold899/A sky130_fd_sc_hd__mux2_1
XANTENNA_fanout151_X fanout151/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_X fanout249/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout530_A fanout538/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_A2 fanout478/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[11\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[15\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1164/X m_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout585/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout416_X fanout416/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout282/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_37_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold777/X fanout205/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_1135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1125/A fanout65/X fanout77/X hold558/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout64_X fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold427/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_701 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__and3_2_B m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__a22oi_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[39\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[40\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_1
XFILLER_56_881 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_43_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__a211oi_2_C1
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y/A1
+ fanout105/X ANTENNA_3/DIODE m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_71_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_350 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X
+ fanout187/X m_blake2.m_hash256.h_flat\[161\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[225\]_sky130_fd_sc_hd__nand2_2_B/Y
+ fanout274/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ sky130_fd_sc_hd__o2bb2a_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y
+ hold933/A fanout84/X fanout144/X m_blake2.m_hash256.m_matrix\[10\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X/A1
+ sky130_fd_sc_hd__a221oi_1
XFILLER_16_778 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X
+ m_blake2.m_hash256.m_g.a0\[20\]_sky130_fd_sc_hd__xor2_2_X/B m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y/A2
+ m_blake2.m_hash256.m_g.a0\[23\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[24\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_11_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold135/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1018/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold429/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_465 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_988 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
XFILLER_48_1013 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold192/X fanout319/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[186\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout190/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B fanout487/X m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_38_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold758/A fanout108/X fanout120/X m_blake2.m_hash256.m_matrix\[15\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_4_1140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1226/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__a22o_2_A1 hold473/A fanout291/X
+ fanout285/X hold449/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_80_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.res_cnt_q\[0\]_sky130_fd_sc_hd__xor2_2_B fanout446/X m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C/B
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__xor2_1
XFILLER_59_1153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__nor2_2_B_A fanout500/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[12\]\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold636/X fanout226/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1_A1
+ m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0 hold455/A m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__mux2_1_A1/X
+ fanout372/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__and3_2_C_A fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X/A
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X/B
+ m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1/A2
+ sky130_fd_sc_hd__or3_2
Xhold922 hold922/A VGND VGND VPWR VPWR hold922/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout209_A fanout212/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout111_A fanout111/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold911 hold911/A VGND VGND VPWR VPWR hold911/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold900 hold900/A VGND VGND VPWR VPWR hold900/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 hold944/A VGND VGND VPWR VPWR hold944/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 hold955/A VGND VGND VPWR VPWR hold955/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[1\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1192/X hold1133/X fanout554/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold43/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xhold933 hold933/A VGND VGND VPWR VPWR hold933/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[14\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold973/A sky130_fd_sc_hd__dfxtp_1
Xhold977 hold977/A VGND VGND VPWR VPWR hold977/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold988 hold988/A VGND VGND VPWR VPWR hold988/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__mux2_1_A0 hold273/A m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold966 hold966/A VGND VGND VPWR VPWR hold966/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[10\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold1137/X m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout235/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_44_1400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold999 hold999/A VGND VGND VPWR VPWR hold999/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout480_A fanout480/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1062 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold441/X m_blake2.m_hash256.v_q\[3\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout416/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_56_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_C1
+ fanout354/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__mux2_1_A0 hold162/X hold852/A
+ fanout571/X VGND VGND VPWR VPWR hold163/A sky130_fd_sc_hd__mux2_1
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__a22o_2_A1 hold548/A fanout192/X
+ fanout198/X hold587/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout24_A fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold564/X fanout563/X
+ VGND VGND VPWR VPWR hold565/A sky130_fd_sc_hd__mux2_1
XFILLER_12_214 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[10\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[10\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1236/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__and3_2_C_A fanout447/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_1437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__mux2_1_A0 hold295/X m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_10_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__xor2_2_B hold1127/A hold498/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.g_buffer\[4\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_49_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold940/X m_blake2.m_hash256.v_q\[15\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[12\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[11\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.v_q\[11\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold430/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold568/A m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout396/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_S fanout414/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold333/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1046/X fanout220/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B fanout484/X hold229/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[5\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
XFILLER_15_1023 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_8_763 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[5\]\[21\]_sky130_fd_sc_hd__xor2_2_A/B sky130_fd_sc_hd__dfxtp_1
Xhold207 hold207/A VGND VGND VPWR VPWR hold207/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__mux2_1_A1_S fanout330/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold218 hold218/A VGND VGND VPWR VPWR hold218/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__a22o_2_B2 hold1245/A fanout265/X fanout305/X
+ m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__a22o_2_B2/X
+ sky130_fd_sc_hd__a22o_1
Xhold229 hold229/A VGND VGND VPWR VPWR hold229/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold242/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold612/X fanout206/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[1\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold885/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.v_q\[12\]\[11\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D
+ fanout424/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a311o_2_B1
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[18\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__a21o_2_X/A2
+ sky130_fd_sc_hd__a311o_1
XFILLER_61_1043 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold949/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[15\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold263/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold927/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.v_q\[4\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold209/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout159_A fanout160/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.h_flat\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold130/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold824/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout182/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_79_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_1145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_fanout326_A fanout342/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold836/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1
+ fanout268/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold207/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout114_X fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout1 fanout1/A VGND VGND VPWR VPWR fanout1/X sky130_fd_sc_hd__buf_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_S fanout211/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold730 hold730/A VGND VGND VPWR VPWR hold730/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 hold741/A VGND VGND VPWR VPWR hold741/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold752 hold752/A VGND VGND VPWR VPWR hold752/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[11\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold421/X hold613/A fanout563/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold763 hold763/A VGND VGND VPWR VPWR hold763/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold774 hold774/A VGND VGND VPWR VPWR hold774/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 hold796/A VGND VGND VPWR VPWR hold796/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1 sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1079/X hold900/X fanout555/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold785 hold785/A VGND VGND VPWR VPWR hold785/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_76_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[30\]_sky130_fd_sc_hd__xor2_2_X/A
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold887/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[181\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__xnor2_2_A hold356/A hold879/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.g_buffer\[12\].m_c_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_79_1337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__mux2_1_A0 hold45/A m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[227\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_73_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3
+ fanout469/X fanout474/X m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout345/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
Xm_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[11\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_4_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout420/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout295/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__mux2_1_A0 hold69/A m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout504/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[127\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_68_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__or2_2_B fanout494/X hold157/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[101\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_71_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[24\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout181/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout27_X fanout27/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1078 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_1067 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or3_2_C
+ fanout346/X m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/A2
+ sky130_fd_sc_hd__or3_1
XFILLER_13_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[7\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1056/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold930/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_1267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__a21o_2_B1 m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/C m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_C1
+ fanout178/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold85/A sky130_fd_sc_hd__dfxtp_1
Xhold90 hold90/A VGND VGND VPWR VPWR hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold424/X hold497/X fanout586/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[9\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold353/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold292/X m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout154/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold88/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout402/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[13\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XFILLER_44_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XFILLER_31_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_14_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1 m_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1/X m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold744/A fanout52/X fanout32/X hold784/A m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout258/X m_blake2.m_hash256.v_q\[6\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout381/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[31\]_sky130_fd_sc_hd__mux2_1_A1_S fanout224/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[12\].m_c_buf m_blake2.m_hash256.g_buffer\[12\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[12\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_67_1241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D_sky130_fd_sc_hd__o31a_2_X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/C m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/D
+ sky130_fd_sc_hd__o31a_1
Xm_blake2.m_hash256.m_matrix\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1200/X m_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout580/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_70_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout506 fanout507/X VGND VGND VPWR VPWR fanout506/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__and3_2_A_B fanout465/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout539 fanout539/A VGND VGND VPWR VPWR fanout539/X sky130_fd_sc_hd__buf_4
XFILLER_59_707 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout528 fanout529/X VGND VGND VPWR VPWR fanout528/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__xor2_4
Xfanout517 fanout519/X VGND VGND VPWR VPWR fanout517/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout201/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B
+ fanout408/X fanout249/X VGND VGND VPWR VPWR fanout173/A sky130_fd_sc_hd__nor2_2
Xm_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__o21a_2_X
+ hold816/A fanout381/X fanout193/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__o21a_1
XFILLER_67_762 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout276_A fanout276/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_S fanout231/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A0 hold110/A m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout518/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold803/A fanout28/X fanout36/X hold918/A m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_16_Left_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_25_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold817/A fanout32/X fanout40/X hold771/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_22_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout610_A fanout615/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__a22o_2_A1/B1 sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_d\[5\]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout186/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout231_X fanout231/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__or4_2
Xm_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
Xm_blake2.m_hash256.m_matrix\[10\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold630/X m_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout578/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold518/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold220/X fanout165/X m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[39\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xhold560 hold560/A VGND VGND VPWR VPWR hold560/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold571 hold571/A VGND VGND VPWR VPWR hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 hold593/A VGND VGND VPWR VPWR hold593/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold582 hold582/A VGND VGND VPWR VPWR hold582/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B fanout486/X hold258/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1136/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2_A1 m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1260 hold1260/A VGND VGND VPWR VPWR hold1260/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1093 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.c_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout24/X fanout52/X
+ hold962/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout132/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_3_X_sky130_fd_sc_hd__o31a_2_A3
+ fanout453/X fanout455/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_3/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y
+ fanout160/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_A1
+ fanout267/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_75_1009 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_695 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y
+ hold603/A fanout377/X fanout185/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/A1
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[15\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__o211a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_A2 m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B
+ fanout402/X m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[41\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1/C1
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[12\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout192/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_S fanout154/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[19\]_sky130_fd_sc_hd__and4_2_C/C
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_1280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_710 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_S fanout159/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_blake2.m_hash256.h_flat\[11\]_sky130_fd_sc_hd__o22a_2_A2/X
+ hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout320/X VGND VGND VPWR VPWR hash\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[15\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold549/X data\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout560/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_matrix\[15\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__mux2_1
XFILLER_17_681 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold601/A fanout110/X fanout94/X hold926/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_20_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1 m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/A2
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/X
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0 hold813/X m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout299/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1
+ m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__a211o_2_A1/X m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout404/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_2
XFILLER_69_1325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__a221o_2_A1 hold464/A fanout289/X
+ fanout277/X hold734/A m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__and3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_30_1137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout412/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1253/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__a22o_2_B2_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
XANTENNA_m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2
+ fanout168/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold536/X fanout587/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout314 fanout342/A VGND VGND VPWR VPWR fanout314/X sky130_fd_sc_hd__buf_2
Xfanout303 fanout303/A VGND VGND VPWR VPWR fanout303/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.h_flat\[253\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold713/A sky130_fd_sc_hd__dfxtp_1
Xfanout336 fanout341/X VGND VGND VPWR VPWR fanout336/X sky130_fd_sc_hd__buf_4
Xfanout347 fanout349/X VGND VGND VPWR VPWR fanout347/X sky130_fd_sc_hd__buf_2
XANTENNA_fanout393_A fanout398/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__or2_2_B_A fanout492/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_1127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout325 fanout326/X VGND VGND VPWR VPWR fanout325/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B sky130_fd_sc_hd__dfxtp_2
Xfanout369 fanout370/X VGND VGND VPWR VPWR fanout369/X sky130_fd_sc_hd__buf_2
Xfanout358 fanout361/X VGND VGND VPWR VPWR fanout358/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout181_X fanout181/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout195/X m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[177\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout187/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout279_X fanout279/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_968 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1/B1 m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_905 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout446_X fanout446/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_735 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__and3_2_C fanout447/X fanout480/X
+ hold165/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X
+ fanout107/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_1173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold923/A fanout109/X fanout88/X m_blake2.m_hash256.m_matrix\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_971 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_46_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nor2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/Y m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[4\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2/A1
+ sky130_fd_sc_hd__nor2_1
XFILLER_7_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_buffer\[13\].m_y_buf m_blake2.m_hash256.g_buffer\[13\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[13\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xm_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__or2_2_A/A fanout162/X m_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout614/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_52_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__mux2_1_A0_S fanout234/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold390 hold390/A VGND VGND VPWR VPWR hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_1111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout94_X fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__mux2_1_A1 hold130/A m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout489/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold999/X m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout155/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/A
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A/X m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/Y
+ sky130_fd_sc_hd__nor3_1
Xm_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B fanout429/X hold249/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout175/X hold787/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[15\].m_c_buf/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_19_946 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ hold401/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_46_776 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1090 hold1090/A VGND VGND VPWR VPWR hold1090/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_73_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout69/X fanout73/X
+ hold984/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__xnor2_2_A hold322/A hold731/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1196/X m_blake2.m_hash256.m_matrix\[10\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout544/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_20_clk_A clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1197/A fanout31/X fanout71/X m_blake2.m_hash256.m_matrix\[7\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold82/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__and3_2_A hold359/A fanout463/X fanout368/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__a211oi_2_A1_C1 fanout371/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C/A
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold428/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[167\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold651/X fanout338/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[159\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_1364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[210\]_sky130_fd_sc_hd__and2_2_B_A fanout432/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X m_blake2.m_hash256.h_flat\[71\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1204/X m_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout568/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
XFILLER_7_1193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B fanout499/X m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold122/X fanout313/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_58_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_25_949 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold351/X m_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout560/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B/A
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A/B sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A1_S fanout411/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout239_A fanout239/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/C
+ m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/B
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_3
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR fanout139/A sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_41_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__a21oi_2_B1/Y VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[3\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
XANTENNA_fanout406_A fanout406/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_c_buf\[2\]_sky130_fd_sc_hd__a211o_2_X m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ m_blake2.m_hash256.g_c_buf\[2\]_sky130_fd_sc_hd__a211o_2_X/A2 m_blake2.m_hash256.v_q\[8\]\[2\]_sky130_fd_sc_hd__o21a_2_A1/X
+ m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__o21a_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[2\].m_c_buf/A sky130_fd_sc_hd__a211o_1
Xm_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor2_2_Y m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/X
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B VGND
+ VGND VPWR VPWR m_io.m_config.nn_q\[3\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold1096/A fanout138/X fanout150/X m_blake2.m_hash256.m_matrix\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A0 hold94/A m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_54_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__o211a_2_C1
+ fanout449/X m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C
+ m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1/C1
+ sky130_fd_sc_hd__o211a_1
XFILLER_47_1420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout122 fanout123/X VGND VGND VPWR VPWR fanout122/X sky130_fd_sc_hd__clkbuf_4
Xfanout111 fanout111/A VGND VGND VPWR VPWR fanout111/X sky130_fd_sc_hd__clkbuf_2
Xfanout100 fanout103/X VGND VGND VPWR VPWR fanout100/X sky130_fd_sc_hd__buf_6
XFILLER_75_805 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout138/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold1047/X fanout308/X VGND VGND VPWR VPWR data\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout144 fanout147/A VGND VGND VPWR VPWR fanout144/X sky130_fd_sc_hd__buf_4
Xfanout133 fanout135/A VGND VGND VPWR VPWR fanout133/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.m_matrix\[7\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold780/X hold1073/A fanout571/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout155 fanout156/X VGND VGND VPWR VPWR fanout155/X sky130_fd_sc_hd__buf_4
XFILLER_75_816 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout166 fanout167/X VGND VGND VPWR VPWR fanout166/X sky130_fd_sc_hd__buf_2
Xfanout199 fanout200/X VGND VGND VPWR VPWR fanout199/X sky130_fd_sc_hd__clkbuf_4
Xfanout177 fanout180/A VGND VGND VPWR VPWR fanout177/X sky130_fd_sc_hd__buf_4
Xfanout188 fanout189/X VGND VGND VPWR VPWR fanout188/X sky130_fd_sc_hd__clkbuf_4
Xm_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__or2_2_A hold307/A fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[32\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_41_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B fanout483/X hold75/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[81\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_c_buf\[11\]_sky130_fd_sc_hd__a221o_2_X hold726/A fanout174/X
+ m_blake2.m_hash256.g_c_buf\[25\]_sky130_fd_sc_hd__a22o_2_X/A2 hold695/A m_blake2.m_hash256.g_c_buf\[11\]_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[11\].m_c_buf/A sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__or2_2_B_A fanout485/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2 m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/A1
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/A2 m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/A3
+ fanout100/X hold459/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/X
+ sky130_fd_sc_hd__o32a_2
XFILLER_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_993 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold871/A fanout116/X fanout96/X hold513/A m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ fanout198/X m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout190/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_13_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__nor2_1
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[97\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold80/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout183/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold115/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[98\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__a22o_2_A1 hold557/A fanout293/X
+ fanout287/X hold692/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_78_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold626/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B/A
+ hold340/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_77_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_1 fanout462/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o21a_2_A1_1/X sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.b_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/B
+ m_blake2.m_hash256.m_g.c_q\[10\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XFILLER_61_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/A
+ m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__nor3b_2_C_N/B m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__nor3b_1
Xm_blake2.m_hash256.m_matrix\[15\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold814/X data\[3\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout559/X VGND VGND VPWR VPWR
+ hold815/A sky130_fd_sc_hd__mux2_1
XFILLER_34_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout353/X m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__a22o_2_A1/X fanout180/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[118\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[126\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y/A m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__a22o_2_A1 hold419/A fanout187/X
+ fanout195/X hold796/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[4\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout307/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__a211o_2_A1 hold496/A fanout280/X
+ m_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__a22o_2_A1/X fanout389/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[3\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[95\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[103\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_57_827 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout189_A fanout192/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout91/X fanout99/X
+ hold1111/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y
+ fanout512/X m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[130\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ sky130_fd_sc_hd__nand2_1
XANTENNA_hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_Q hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A fanout361/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_buffer\[13\].m_y_buf/A sky130_fd_sc_hd__o32a_1
XANTENNA_fanout523_A fanout524/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_738 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_X fanout144/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold762/X fanout555/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_1441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout409_X fanout409/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_5_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload3/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1232/A sky130_fd_sc_hd__dfxtp_1
Xm_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.cmd\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold1236/A fanout145/X fanout97/X hold1243/A m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[65\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[73\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/B sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_0_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_1147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ hold917/A fanout137/X fanout121/X hold1006/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_74_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold748/A fanout29/X fanout77/X hold889/A m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[6\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_47_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XFILLER_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout106/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold843/X m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_4_Left_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_941 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_1118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 hold715/X m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout302/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout24/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1 hold738/A fanout349/X
+ fanout260/X m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1/B2 fanout268/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1170/X
+ fanout586/X VGND VGND VPWR VPWR hold1171/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR fanout51/A sky130_fd_sc_hd__nor2_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_S fanout155/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_1269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0 hold740/X m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout417/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_1016 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__o21ai_2_A1_B1 fanout193/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.v_q\[0\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold878/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
XFILLER_62_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_34_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ hold1131/A fanout78/X m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout22/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XFILLER_37_1452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold455/X fanout410/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_matrix\[11\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[11\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold522/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout221/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold47/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold892/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold432/X m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold912 hold912/A VGND VGND VPWR VPWR hold912/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold901 hold901/A VGND VGND VPWR VPWR hold901/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold945 hold945/A VGND VGND VPWR VPWR hold945/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout104_A fanout107/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold923 hold923/A VGND VGND VPWR VPWR hold923/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 hold934/A VGND VGND VPWR VPWR hold934/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 hold978/A VGND VGND VPWR VPWR hold978/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold967 hold967/A VGND VGND VPWR VPWR hold967/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 hold956/A VGND VGND VPWR VPWR hold956/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold989 hold989/A VGND VGND VPWR VPWR hold989/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold663/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__nand2_2_B fanout440/X hold230/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[183\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_44_1412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C
+ m_blake2.m_hash256.m_g.c_q\[30\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C/B
+ m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/B sky130_fd_sc_hd__nand3_2
Xm_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1/B1
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__o211a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout109/X
+ fanout149/X hold1223/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_32_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1052 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_32_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_32_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold532/X m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout299/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1036/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR
+ VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__dfxtp_1
XFILLER_53_841 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold92/A m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout504/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_77_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_A_N m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_A_N/X sky130_fd_sc_hd__and2b_1
XANTENNA_m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.h_flat\[132\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold221/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold858/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_709 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ hold910/X VGND VGND VPWR VPWR hold909/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__and3_2_C_B fanout480/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[68\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout25/X fanout69/X
+ hold923/A m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_23_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[15\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ data\[4\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR data\[4\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o21a_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1/B1
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_5_926 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.v_q\[14\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold664/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold1129/X m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout156/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__and2b_2_B_A_N
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[2\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold472/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2
+ fanout266/X m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[60\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout267/A VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[92\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[22\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A
+ m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1 hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[19\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[29\]_sky130_fd_sc_hd__or2_2_A hold303/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[29\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold568/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold149/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold164/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[201\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2_A2 fanout265/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[4\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1094/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_720 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[8\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[15\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold787/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__mux2_1_A0 hold301/X m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout231/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[13\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold497/X hold786/X fanout582/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold328/A fanout36/X fanout44/X hold920/A m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold208 hold208/A VGND VGND VPWR VPWR hold208/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[8\]\[16\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1203/X fanout221/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold219 hold219/A VGND VGND VPWR VPWR hold219/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout213/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_1309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold771/X hold515/X fanout554/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_28_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__and2_2_B fanout439/X hold94/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[14\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold538/X m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout210/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_39_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[12\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_79_793 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout478/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold929/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.d_q\[6\]_sky130_fd_sc_hd__xor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold296/A m_blake2.m_hash256.h_flat\[213\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout397/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_67_999 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__nor2_2_B_A fanout484/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__inv_2_Y fanout606/X
+ VGND VGND VPWR VPWR m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X/B1 sky130_fd_sc_hd__inv_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout302/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_830 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload21/A m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__a32o_2_A1_A2 fanout354/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[13\]_sky130_fd_sc_hd__o22a_2_A2/B1
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold954/X hold729/X fanout600/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/A
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/B
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_20_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1 hold679/A fanout377/X
+ fanout193/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2_sky130_fd_sc_hd__o21bai_2_Y_Y
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A fanout222/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[31\]_sky130_fd_sc_hd__xor2_2_B/X
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[14\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold939/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_buffer\[0\].m_c_buf m_blake2.m_hash256.g_buffer\[0\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[0\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[8\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold983/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X
+ fanout194/X m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout186/X fanout273/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1 m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ fanout451/X m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1/X
+ sky130_fd_sc_hd__o31a_1
Xhold720 hold720/A VGND VGND VPWR VPWR hold720/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__and3_2_B hold1254/A
+ m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1 m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__and2_2_A/B
+ sky130_fd_sc_hd__and3_1
Xhold731 hold731/A VGND VGND VPWR VPWR hold731/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 hold753/A VGND VGND VPWR VPWR hold753/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 hold764/A VGND VGND VPWR VPWR hold764/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold742 hold742/A VGND VGND VPWR VPWR hold742/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 hold797/A VGND VGND VPWR VPWR hold797/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout590_A fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold786 hold786/A VGND VGND VPWR VPWR hold786/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 hold775/A VGND VGND VPWR VPWR hold775/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.h_flat\[226\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold73/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__and2_2_B_A fanout430/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2 m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ fanout265/X fanout305/X hold642/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_fanout476_X fanout476/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[105\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold290/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[235\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0_S
+ fanout520/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_969 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/Y sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_68_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[114\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold69/X fanout311/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_874 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout402/X m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__a211o_2_A1/X
+ m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A2_N
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_64_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a221o_2_C1
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a221o_2_C1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[7\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[9\]_sky130_fd_sc_hd__a211oi_2_A1_A2 fanout402/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__nor3_2_Y
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__nor3_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1_sky130_fd_sc_hd__a21o_2_A2/B1
+ sky130_fd_sc_hd__nand2_1
XFILLER_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/B m_blake2.m_hash256.m_g.a_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.g_c_buf\[6\]_sky130_fd_sc_hd__a211o_2_X_A1 m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.c_q\[14\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/B
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A/C sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout126/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[5\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/A1 m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1196/A fanout32/X fanout76/X hold1123/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_955 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[8\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1123/X hold1165/A fanout551/X VGND VGND VPWR VPWR hold1124/A sky130_fd_sc_hd__mux2_1
XFILLER_76_774 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold91 hold91/A VGND VGND VPWR VPWR hold91/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A0 hold87/A m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout508/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_io.m_config.ll_q\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X hold1106/X
+ VGND VGND VPWR VPWR hold505/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold80 hold80/A VGND VGND VPWR VPWR hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A0 hold960/A m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__xnor2_2_A hold439/A hold1150/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_1_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout360/X m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a21o_1
XFILLER_50_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_833 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout284/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_70_clk clkload0/A VGND VGND VPWR VPWR clkload12/A sky130_fd_sc_hd__clkbuf_8
Xm_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2 m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ fanout265/X fanout305/X hold1042/A m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/C1
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/X sky130_fd_sc_hd__a221o_1
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[7\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1073/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X_A2 fanout275/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout507 fanout508/X VGND VGND VPWR VPWR fanout507/X sky130_fd_sc_hd__buf_2
Xfanout529 fanout530/X VGND VGND VPWR VPWR fanout529/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.g_buffer\[16\].m_c_buf m_blake2.m_hash256.g_buffer\[16\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[16\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xfanout518 fanout519/X VGND VGND VPWR VPWR fanout518/X sky130_fd_sc_hd__clkbuf_2
Xm_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__and3_2_A hold1235/A fanout464/X fanout384/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[36\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold530/A fanout42/X fanout78/X hold577/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[26\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold433/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_1033 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[1\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/B2 sky130_fd_sc_hd__o21ai_2
Xm_blake2.m_hash256.m_matrix\[9\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A hold586/X
+ VGND VGND VPWR VPWR hold585/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_1_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout171_A fanout173/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[53\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold110/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[45\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout269_A fanout269/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout182/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/X m_blake2.m_hash256.v_q\[3\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_78_1382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout436_A fanout443/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_1208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_855 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_61_clk clkload2/A VGND VGND VPWR VPWR clkbuf_leaf_61_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B
+ m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.g_buffer\[9\].m_c_buf/X
+ VGND VGND VPWR VPWR ANTENNA_8/DIODE sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout224_X fanout224/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1084/X m_blake2.m_hash256.m_matrix\[6\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout564/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout284/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[174\]_sky130_fd_sc_hd__mux2_1_A1_S fanout328/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A fanout467/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__and2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_C1
+ fanout355/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold238/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_57_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold572 hold572/A VGND VGND VPWR VPWR hold572/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 hold550/A VGND VGND VPWR VPWR hold550/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold561 hold561/A VGND VGND VPWR VPWR hold561/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 hold583/A VGND VGND VPWR VPWR hold583/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 hold594/A VGND VGND VPWR VPWR hold594/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout192/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout200/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout84_A fanout87/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1261 hold1261/A VGND VGND VPWR VPWR hold1261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1250 hold1250/A VGND VGND VPWR VPWR hold1250/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A0 hold43/A m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout529/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_1370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__or2_2_A hold257/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[62\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XFILLER_14_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_buffer\[1\].m_y_buf m_blake2.m_hash256.g_buffer\[1\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[1\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_52_clk clkload3/A VGND VGND VPWR VPWR clkbuf_leaf_52_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__a211oi_2_A1 hold380/A fanout284/X
+ m_blake2.m_hash256.v_q\[1\]\[8\]_sky130_fd_sc_hd__a22o_2_A1/X fanout371/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__a211oi_2_A1/Y sky130_fd_sc_hd__a211oi_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout286/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__a31o_2_B1_A3
+ m_blake2.m_hash256.block_idx_plus_one_q\[43\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_12_1027 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X hold453/A fanout18/X m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X/B2 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[10\].m_y_buf/A sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[23\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[7\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.g_c_buf\[18\]_sky130_fd_sc_hd__a2111o_2_X hold837/A fanout174/X
+ m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.v_q\[11\]\[18\]_sky130_fd_sc_hd__o21a_2_A1/X
+ m_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__o21a_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.g_buffer\[18\].m_c_buf/A sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1186/X
+ fanout587/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1138/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_2
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold893/A fanout140/X fanout116/X m_blake2.m_hash256.m_matrix\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[86\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_48_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_X m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_671 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_19_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold816/A sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_43_clk clkload5/A VGND VGND VPWR VPWR clkbuf_leaf_43_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout268/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_9_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_20_825 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A block_first_sky130_fd_sc_hd__a22o_2_B2/X
+ VGND VGND VPWR VPWR fanout500/A sky130_fd_sc_hd__dfxtp_4
XANTENNA_m_io.m_config.ll_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2
+ fanout163/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a32o_2_X_A1
+ fanout463/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.fsm_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a32o_2_X_B2
+ fanout478/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[203\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[6\]\[3\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout520/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[12\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__or2_2_A hold490/A fanout376/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_d\[13\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1
+ fanout269/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__xnor2_2_A hold592/A hold777/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.g_buffer\[15\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold211/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__a31o_2_A3 fanout448/X fanout479/X
+ hold208/A fanout512/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_A m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout275/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout304 fanout307/A VGND VGND VPWR VPWR fanout304/X sky130_fd_sc_hd__clkbuf_4
XFILLER_67_1061 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A0 hold89/A m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout518/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xfanout315 fanout316/X VGND VGND VPWR VPWR fanout315/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__xnor2_2_A hold507/A hold1262/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xfanout348 fanout349/X VGND VGND VPWR VPWR fanout348/X sky130_fd_sc_hd__clkbuf_2
Xfanout337 fanout338/X VGND VGND VPWR VPWR fanout337/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout326 fanout342/X VGND VGND VPWR VPWR fanout326/X sky130_fd_sc_hd__buf_2
Xfanout359 fanout361/X VGND VGND VPWR VPWR fanout359/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload31/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__a22o_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_52_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[2\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1134/X hold1270/X fanout553/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_C1
+ fanout177/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_914 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout174_X fanout174/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__and2_2_B fanout442/X hold59/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[22\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_55_799 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__o21ai_2_Y
+ fanout469/X m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ fanout481/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y/B1
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout341_X fanout341/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_34_clk clkload4/A VGND VGND VPWR VPWR clkbuf_leaf_34_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_4
XFILLER_74_1087 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B/Y m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__xnor2_2_A hold836/A hold1098/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout18/X hold1004/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[16\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA_m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1_A2
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_46_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold856/X fanout541/X
+ VGND VGND VPWR VPWR hold857/A sky130_fd_sc_hd__mux2_1
XFILLER_10_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_59_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__xor2_2_A hold859/A hold260/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_59_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[0\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_buffer\[17\].m_y_buf m_blake2.m_hash256.g_buffer\[17\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[17\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.g_b\[0\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1222/X hold1211/X fanout580/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold380 hold380/A VGND VGND VPWR VPWR hold380/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold391 hold391/A VGND VGND VPWR VPWR hold391/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_A fanout486/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout52/X
+ fanout76/X hold1136/A m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__xnor2_2_A hold904/A hold501/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__nor2_2_B fanout492/X hold169/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[228\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_2
Xhold1080 hold1080/A VGND VGND VPWR VPWR hold1080/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1091 hold1091/A VGND VGND VPWR VPWR hold1091/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_4
XTAP_TAPCELL_ROW_16_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clkload1/A VGND VGND VPWR VPWR clkbuf_leaf_25_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_61_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold621/X fanout585/X
+ VGND VGND VPWR VPWR hold622/A sky130_fd_sc_hd__mux2_1
XFILLER_14_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout198/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_663 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y m_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a0\[21\]_sky130_fd_sc_hd__xnor2_2_Y/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold729/A fanout58/X fanout27/X hold757/A m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_862 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X
+ fanout1/X fanout610/X input5/X VGND VGND VPWR VPWR m_io.m_config.data_i\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__a22o_2_A1/B1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_6_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/B m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y
+ sky130_fd_sc_hd__nand3b_4
XPHY_EDGE_ROW_79_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_869 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_847 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold360/X fanout168/X m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__or2_2_A/X fanout620/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__nor2_2_B_A fanout499/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_722 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout153/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout28/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout200/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[3\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout56/X m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a2111o_1
XFILLER_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold988/A fanout86/X fanout90/X hold1058/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_16_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_16_clk/X sky130_fd_sc_hd__clkbuf_8
XFILLER_51_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR fanout135/A sky130_fd_sc_hd__and4_2
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_2
XTAP_TAPCELL_ROW_41_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1082 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_1071 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B fanout408/X hold598/A
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/X sky130_fd_sc_hd__and3_1
XFILLER_20_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.h_flat\[164\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold53/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout301_A fanout303/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__a31o_2_B1_B1
+ m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_54_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/C
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__and2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1/B1 sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold680/A fanout33/X fanout41/X m_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[15\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold94/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[165\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xfanout101 fanout103/X VGND VGND VPWR VPWR fanout101/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xfanout112 fanout115/A VGND VGND VPWR VPWR fanout112/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0/X
+ m_blake2.m_hash256.v_q\[0\]\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.h_flat\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1 sky130_fd_sc_hd__xnor2_1
Xfanout123 fanout123/A VGND VGND VPWR VPWR fanout123/X sky130_fd_sc_hd__buf_2
XFILLER_59_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout134 fanout135/A VGND VGND VPWR VPWR fanout134/X sky130_fd_sc_hd__clkbuf_4
Xfanout145 fanout147/A VGND VGND VPWR VPWR fanout145/X sky130_fd_sc_hd__buf_2
XANTENNA_fanout291_X fanout291/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout156 fanout156/A VGND VGND VPWR VPWR fanout156/X sky130_fd_sc_hd__buf_4
Xm_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[7\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold495/A sky130_fd_sc_hd__dfxtp_1
Xfanout167 fanout168/X VGND VGND VPWR VPWR fanout167/X sky130_fd_sc_hd__buf_2
Xfanout189 fanout192/A VGND VGND VPWR VPWR fanout189/X sky130_fd_sc_hd__clkbuf_4
Xfanout178 fanout180/A VGND VGND VPWR VPWR fanout178/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_1031 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_744 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__mux2_1_A0_S fanout301/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_906 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout47_A fanout47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout60/X m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout20/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_48_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1225/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X
+ fanout87/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_666 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__or2_2_A hold575/A fanout387/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[30\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_13_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B fanout206/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XFILLER_3_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_A1
+ fanout278/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__and2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout140/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__a21oi_2
Xm_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout241/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_2_1091 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[10\]_sky130_fd_sc_hd__or2_2_A hold317/A fanout242/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[10\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout201/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1250/X
+ fanout554/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__nand2b_2_B m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_1
Xm_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A hold877/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__mux2_1_A1_S fanout215/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__xor2_2_A hold755/A hold874/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout414/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkload7/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__a22o_2_A1 hold367/A fanout290/X
+ fanout284/X hold431/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR uo_out[7] sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1
+ fanout348/X m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2/X
+ m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X fanout255/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ sky130_fd_sc_hd__a2bb2o_1
Xm_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ hold555/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__or2_2_A hold760/A fanout372/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[12\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_68_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1097 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/D m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold811/X hold970/A fanout573/X VGND VGND VPWR VPWR hold812/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout416/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_71_clk/X
+ m_blake2.m_hash256.m_matrix\[8\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold889/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0 hold279/A m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout362/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[153\]_sky130_fd_sc_hd__and2_2_B_A fanout430/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1237/X m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_B
+ fanout445/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3/B1 VGND VGND
+ VPWR VPWR fanout184/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout251_A fanout252/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout349_A fanout350/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_43_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__mux2_1_A0 hold17/A m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout536/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout516_A fanout539/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold323/X m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout236/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_1453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[20\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[38\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout114/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__mux2_1_A0 hold1014/X m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout413/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_1328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A_B m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1 m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/B1
+ m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/B2 m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__o211a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1/Y
+ sky130_fd_sc_hd__a221oi_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__and3_2_B m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/A1
+ m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__a2bb2o_2_A1_N/B2 m_blake2.m_hash256.block_idx_plus_one_q\[54\]_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/C
+ sky130_fd_sc_hd__and3_1
XFILLER_48_806 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__a22o_2_A1 hold440/A fanout189/X
+ fanout197/X hold610/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X
+ fanout99/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_1159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1041/X m_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout569/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__xor2_2_B hold996/A hold496/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[15\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[10\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold629/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_1446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout102/X hold683/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__o32a_2
XFILLER_16_725 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__mux2_1_A0 hold251/X m_blake2.m_hash256.v_q\[7\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout230/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold361/A fanout92/X fanout148/X hold1113/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[5\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__a21o_2_B1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/C sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.d_q\[7\]_sky130_fd_sc_hd__xor2_2_B/X m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout184/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_34_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_A2 fanout289/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold501/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_913 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.g_buffer\[9\].m_y_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[9\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XANTENNA_clkbuf_leaf_49_clk_A clkload2/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[7\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1208/X hold1266/A fanout544/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1_S fanout202/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ hold494/X VGND VGND VPWR VPWR hold493/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[14\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.v_q\[11\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1100/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1062/X fanout217/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold616/A sky130_fd_sc_hd__dfxtp_1
XFILLER_78_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_S fanout419/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_669 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_2
Xm_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X/A
+ m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold336/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A0 hold191/A m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1006 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold942/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout181/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_864 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold620/A fanout85/X fanout121/X hold886/A m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/A1
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nand2_1
XFILLER_62_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A1
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XFILLER_21_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2
+ fanout267/X m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[79\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2/X
+ fanout389/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[47\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2/Y
+ sky130_fd_sc_hd__o211ai_1
Xm_blake2.m_hash256.v_q\[13\]\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1024/X fanout208/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[1\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[1\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold193/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[16\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold756/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold1036/A fanout30/X fanout75/X hold536/A m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[9\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_2
XFILLER_30_761 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__mux2_1_A0 hold618/X m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout303/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[19\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xhold902 hold902/A VGND VGND VPWR VPWR hold902/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 hold913/A VGND VGND VPWR VPWR hold913/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A1_S fanout327/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__or2_2_B fanout499/X hold82/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1107/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_77_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold924 hold924/A VGND VGND VPWR VPWR hold924/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__and3_2_A/A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A/B VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[7\]_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xhold946 hold946/A VGND VGND VPWR VPWR hold946/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold935 hold935/A VGND VGND VPWR VPWR hold935/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 hold968/A VGND VGND VPWR VPWR hold968/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold979 hold979/A VGND VGND VPWR VPWR hold979/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 hold957/A VGND VGND VPWR VPWR hold957/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhash\[6\]_sky130_fd_sc_hd__or2_2_B fanout500/X hash\[6\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR hash\[6\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold560/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold1127/X fanout219/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[6\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_69_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y/A
+ m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[8\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout299_A fanout299/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold210/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold860/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[3\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold954/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_A1
+ fanout283/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0 hold596/X m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_72_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_861 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkload10/A m_blake2.m_hash256.m_g.a0\[16\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[16\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.m_matrix\[5\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1070/X hold1020/X fanout570/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold92/X fanout312/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.fsm_q\[0\]_sky130_fd_sc_hd__or2_2_B fanout478/X hold185/A VGND
+ VGND VPWR VPWR fanout422/A sky130_fd_sc_hd__or2_4
Xm_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold567/X fanout204/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_52_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout254_X fanout254/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_706 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_80_683 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout421_X fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__a22o_2_A1 hold956/A fanout258/X
+ fanout199/X hold712/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X/A
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND
+ VPWR VPWR hold1261/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X/A2
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout101/X m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/B2 VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ sky130_fd_sc_hd__o32a_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_23_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__xor2_2_B hold640/A hold527/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold374/X m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout159/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[9\]\[18\]_sky130_fd_sc_hd__xor2_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_938 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.g_buffer\[17\].m_c_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.ll_q\[61\]_sky130_fd_sc_hd__and3_2_A_B fanout465/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[11\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold706/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[10\]\[13\]_sky130_fd_sc_hd__o21a_2_A1 hold742/A fanout378/X
+ fanout169/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[13\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__o21a_1
XFILLER_79_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ fanout450/X fanout457/X fanout462/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B fanout486/X hold122/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[13\]\[24\]_sky130_fd_sc_hd__a2bb2o_2_A1_N hold285/A fanout380/X
+ fanout264/X hold1254/A VGND VGND VPWR VPWR m_io.m_config.ll_q\[56\]_sky130_fd_sc_hd__a211o_2_A1/B1
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_48_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_S fanout232/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X
+ hold1074/A fanout90/X fanout138/X hold1133/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout284/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X
+ m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B/B
+ m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout501/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_16_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X hold660/X fanout275/X m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X/C1 VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[1\]_sky130_fd_sc_hd__a211o_2_X/X
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_16_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[12\]\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1210/X fanout227/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.m_matrix\[0\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ hold895/X VGND VGND VPWR VPWR hold894/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ hold243/A fanout305/X m_blake2.m_hash256.v_q\[12\]\[27\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.m_matrix\[13\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1029/X hold1036/A fanout559/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__a211o_2_A1 hold556/A fanout289/X
+ m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__a22o_2_A1/X fanout362/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[16\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XFILLER_67_1424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold209 hold209/A VGND VGND VPWR VPWR hold209/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[14\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold383/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[15\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/D
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X
+ fanout351/X m_blake2.m_hash256.v_q\[5\]\[20\]_sky130_fd_sc_hd__a22o_2_A1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__and2_1
XANTENNA_block_last_sky130_fd_sc_hd__a22o_2_B2_B1_sky130_fd_sc_hd__nor2_2_Y_A fanout422/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ hold912/A fanout54/X fanout78/X hold646/A m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_3_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold463/X m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout153/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold584/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_72_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[2\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A hold1010/X
+ VGND VGND VPWR VPWR hold969/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold296/X fanout215/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__clkinv_2
XFILLER_47_680 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_4_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload2/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__a32o_2_A1_A3 fanout251/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_897 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_50_845 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nor2_2_A/Y m_blake2.m_hash256.m_g.c_q\[17\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A/B
+ sky130_fd_sc_hd__nand2b_1
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[13\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[4\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold620/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[8\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[21\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold597/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold356/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_79_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_79_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_d\[16\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_A2
+ fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_1169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__nor2_2_B fanout484/X hold109/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[104\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_20_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout214_A fanout216/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_1461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[1\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold378/X hold968/A fanout560/X VGND VGND VPWR VPWR hold379/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_11_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold710 hold710/A VGND VGND VPWR VPWR hold710/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[8\]\[22\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold819/X fanout223/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold721 hold721/A VGND VGND VPWR VPWR hold721/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold754 hold754/A VGND VGND VPWR VPWR hold754/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 hold732/A VGND VGND VPWR VPWR hold732/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 hold743/A VGND VGND VPWR VPWR hold743/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_buffer\[4\].m_c_buf m_blake2.m_hash256.g_buffer\[4\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[4\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xhold765 hold765/A VGND VGND VPWR VPWR hold765/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout32/X fanout72/X
+ hold883/A m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout128/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold776 hold776/A VGND VGND VPWR VPWR hold776/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold787 hold787/A VGND VGND VPWR VPWR hold787/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold798 hold798/A VGND VGND VPWR VPWR hold798/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_S fanout156/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_923 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout160/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout371_X fanout371/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_24_Left_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X
+ m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__a221o_2_B2/X
+ m_blake2.m_hash256.v_q\[15\]\[11\]_sky130_fd_sc_hd__o21ai_2_A1/Y fanout268/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_d\[21\]_sky130_fd_sc_hd__nor2_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[21\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_77_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_59_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold791/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold914/A fanout138/X fanout146/X hold1187/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y hash\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_33_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ hold697/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[23\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout424/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[49\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout16/X hold802/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[19\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1_A1 m_blake2.m_hash256.m_g.d_q\[15\]_sky130_fd_sc_hd__xnor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout198/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout90/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_1121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.g_b\[28\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout190/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y/B sky130_fd_sc_hd__a21oi_1
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A m_blake2.m_hash256.h_flat\[232\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold250/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_A1
+ fanout256/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_42_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[25\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2/X
+ m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_C1
+ fanout354/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.h_flat\[111\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold166/A sky130_fd_sc_hd__dfxtp_1
XFILLER_76_786 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[241\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold87/X fanout315/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[233\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[6\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[32\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
Xhold81 hold81/A VGND VGND VPWR VPWR hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A VGND VGND VPWR VPWR hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_1 hold267/A m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout396/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
Xhold92 hold92/A VGND VGND VPWR VPWR hold92/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[13\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[10\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ hold1168/X VGND VGND VPWR VPWR hold1167/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__and2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_c_buf\[18\]_sky130_fd_sc_hd__a2111o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout109/X fanout97/X
+ m_blake2.m_hash256.m_matrix\[6\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[120\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold960/X fanout310/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[112\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2
+ fanout266/X m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.h_flat\[110\]_sky130_fd_sc_hd__nor2_2_B/Y
+ fanout400/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_17_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_992 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X
+ fanout360/X m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X/A2_N
+ m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X fanout257/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X/A1 sky130_fd_sc_hd__a2bb2o_1
XFILLER_17_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_27_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout29/X
+ fanout65/X m_blake2.m_hash256.m_matrix\[11\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[30\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_74_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[3\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__a32o_2_A1_B1 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 ANTENNA_2/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__or2_2_B fanout498/X hold47/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[191\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_28_1205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout508 fanout509/X VGND VGND VPWR VPWR fanout508/X sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_60_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout519 fanout524/X VGND VGND VPWR VPWR fanout519/X sky130_fd_sc_hd__buf_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_1_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__a221o_2_B2_C1 fanout269/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__o21a_2_A1 hold1087/A fanout363/X
+ fanout250/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_1_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout164_A fanout168/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0 hold1190/X m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout296/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[9\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X
+ hold589/A fanout35/X fanout43/X m_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__xnor2_2_A hold455/A hold793/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold574/X m_blake2.m_hash256.m_matrix\[14\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout545/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold988/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__a22o_2_A1 hold775/A fanout174/A
+ m_blake2.m_hash256.v_q\[11\]\[3\]_sky130_fd_sc_hd__or2_2_A/X fanout173/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X/B1 sky130_fd_sc_hd__a22o_1
XANTENNA_fanout429_A fanout431/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout217_X fanout217/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold621/X hold706/X fanout582/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__dfxtp_2_Q clkload19/A m_blake2.m_hash256.h_flat\[137\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold132/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__and3_2_A_X fanout420/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B fanout483/X hold69/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[106\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold540 hold540/A VGND VGND VPWR VPWR hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold562 hold562/A VGND VGND VPWR VPWR hold562/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 hold551/A VGND VGND VPWR VPWR hold551/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 hold584/A VGND VGND VPWR VPWR hold584/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 hold595/A VGND VGND VPWR VPWR hold595/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 hold573/A VGND VGND VPWR VPWR hold573/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[146\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold107/X fanout320/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/A2
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/B1_N
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/Y
+ sky130_fd_sc_hd__o21bai_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_A1
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N/A
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N/Y
+ sky130_fd_sc_hd__nor3b_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold952/A fanout94/X fanout150/X hold732/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold288/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
Xhold1251 hold1251/A VGND VGND VPWR VPWR hold1251/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[13\]_sky130_fd_sc_hd__and4_2_C/A m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2
+ fanout240/X hold364/A m_blake2.m_hash256.v_q\[12\]\[17\]_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[17\]_sky130_fd_sc_hd__a21oi_2_Y/A2 sky130_fd_sc_hd__o221a_1
Xhold1240 hold1240/A VGND VGND VPWR VPWR hold1240/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__a21oi_2_A1/B1 m_blake2.m_hash256.m_g.m_add_1.x2_i\[29\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout108/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xuio_out_sky130_fd_sc_hd__buf_2_X_1 uio_out_sky130_fd_sc_hd__buf_2_X_1/A VGND VGND
+ VPWR VPWR uio_out[7] sky130_fd_sc_hd__buf_2
Xhold1262 hold1262/A VGND VGND VPWR VPWR hold1262/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_73_723 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold43/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[51\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_45_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A1_S fanout409/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout32_X fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__xnor2_2_A hold295/A hold1148/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_buffer\[5\].m_y_buf m_blake2.m_hash256.g_buffer\[5\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[5\].m_y_buf/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X m_io.m_config.ll_q\[43\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1042/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__and2_2_A_A m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A0 hold632/A m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout223/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout186/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[15\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout193/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__xnor2_2_A hold568/A m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[15\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[12\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1122/X hold1152/X fanout552/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X_A2
+ fanout118/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_160 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__xnor2_2_B hold695/A hold318/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_32_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout417/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__and2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_653 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__or2_2_A hold306/A fanout244/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold677/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.res_cnt_q\[0\]_sky130_fd_sc_hd__xor2_2_B_A fanout446/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_1297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[29\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X m_blake2.m_hash256.h_flat\[76\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold280/A sky130_fd_sc_hd__dfxtp_1
XFILLER_69_1349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[1\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold947/X hold757/A fanout573/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/C
+ sky130_fd_sc_hd__and2_1
Xm_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0 m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/Y
+ hold207/A fanout435/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_X_sky130_fd_sc_hd__a31o_2_A3
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1/X
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A1
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout305 fanout307/A VGND VGND VPWR VPWR fanout305/X sky130_fd_sc_hd__clkbuf_2
XFILLER_67_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[85\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold89/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__nand2b_2_A_N_B
+ m_blake2.m_hash256.v_q\[0\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout316 fanout317/X VGND VGND VPWR VPWR fanout316/X sky130_fd_sc_hd__buf_2
Xfanout327 fanout330/X VGND VGND VPWR VPWR fanout327/X sky130_fd_sc_hd__clkbuf_4
Xfanout338 fanout341/X VGND VGND VPWR VPWR fanout338/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.g_buffer\[31\].m_c_buf m_blake2.m_hash256.g_buffer\[31\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[31\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
Xfanout349 fanout350/X VGND VGND VPWR VPWR fanout349/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_52_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X
+ hold934/A fanout108/X m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/B1
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold739/A fanout130/X fanout94/X hold1103/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout281_A fanout282/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A fanout385/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[21\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/A2
+ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout546_A fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.h_flat\[90\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3/X
+ m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[2\]\[26\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[5\]\[15\]_sky130_fd_sc_hd__xor2_2_A/B
+ fanout357/X fanout261/X m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[47\]_sky130_fd_sc_hd__and3_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[15\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__and3_2_B_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[37\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o211a_2_A2
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_B/X
+ fanout468/X fanout401/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A/D
+ sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.v_q\[14\]\[0\]_sky130_fd_sc_hd__mux2_1_A0 hold672/X m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_A_N
+ m_blake2.m_hash256.m_g.b_q\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout289/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_1_clk/X
+ m_blake2.m_hash256.g_buffer\[21\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__a211o_2_A1 hold588/A fanout278/X
+ m_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__a22o_2_A1/X fanout366/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[25\]_sky130_fd_sc_hd__a211o_2_A1/X sky130_fd_sc_hd__a211o_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[4\]_sky130_fd_sc_hd__mux2_1_A1_S fanout207/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__a31o_2_A3 fanout447/X fanout480/X
+ hold171/A fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[142\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[45\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold370 hold370/A VGND VGND VPWR VPWR hold370/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 hold381/A VGND VGND VPWR VPWR hold381/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A0 hold155/A m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout528/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold392 hold392/A VGND VGND VPWR VPWR hold392/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_2_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ hold881/A fanout134/X fanout118/X m_blake2.m_hash256.m_matrix\[13\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2
+ fanout293/X m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2/X
+ fanout356/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[59\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_TAPCELL_ROW_5_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B
+ fanout615/X m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__nand2_2
XFILLER_58_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_block_data.data_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B_sky130_fd_sc_hd__or2_2_X
+ hold4/A m_io.m_block_data.data_cnt_q\[5\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_block_data.data_cnt_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X/B
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2_B1 fanout240/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1092 hold1092/A VGND VGND VPWR VPWR hold1092/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_45_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1070 hold1070/A VGND VGND VPWR VPWR hold1070/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 hold1081/A VGND VGND VPWR VPWR hold1081/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hash\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_Q hash\[6\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[6\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1051/X hold934/X fanout545/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_1190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A/A
+ m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__o211a_2_X
+ hold724/A fanout369/X fanout237/X m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X/C1 sky130_fd_sc_hd__o211a_1
XFILLER_57_1275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_675 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[9\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[11\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_995 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkload7/A m_blake2.m_hash256.m_matrix\[2\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1095/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout300/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_1333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1165/A fanout32/X fanout80/X hold1231/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_69_859 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[9\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold208/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_51_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout102/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X/A
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__o211a_2_X
+ hold809/A fanout381/X fanout239/X m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__a22oi_2_B2/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X/C sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR fanout131/A sky130_fd_sc_hd__and4_2
XANTENNA_fanout127_A fanout127/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[57\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_41_clk/X
+ hold160/X VGND VGND VPWR VPWR hold159/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[4\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1081/X hold1016/X fanout569/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_1381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__or2_2_B fanout492/X hold1189/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[188\]_sky130_fd_sc_hd__or2_2_B/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_54_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_S fanout156/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout102 fanout103/X VGND VGND VPWR VPWR fanout102/X sky130_fd_sc_hd__clkbuf_2
XFILLER_47_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout496_A fanout497/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout113 fanout115/A VGND VGND VPWR VPWR fanout113/X sky130_fd_sc_hd__clkbuf_2
Xm_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout48/X fanout72/X
+ hold933/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[29\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xfanout146 fanout147/A VGND VGND VPWR VPWR fanout146/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_50_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout135 fanout135/A VGND VGND VPWR VPWR fanout135/X sky130_fd_sc_hd__clkbuf_2
Xfanout124 fanout127/A VGND VGND VPWR VPWR fanout124/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_input1_A ena VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout168 fanout168/A VGND VGND VPWR VPWR fanout168/X sky130_fd_sc_hd__buf_2
Xfanout157 fanout160/A VGND VGND VPWR VPWR fanout157/X sky130_fd_sc_hd__buf_4
XFILLER_59_358 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout284_X fanout284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout179 fanout180/X VGND VGND VPWR VPWR fanout179/X sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_35_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_701 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1087 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_48_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_929 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.round_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X
+ fanout456/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/B1
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[19\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold95/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout348/X m_blake2.m_hash256.v_q\[5\]\[26\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ fanout177/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[179\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold145/X fanout322/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout63/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1118/X m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout153/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__xnor2_2_B hold927/A hold704/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[1\]_sky130_fd_sc_hd__xnor2_2_B/Y sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_8_clk_A clkload0/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold609/X fanout587/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__mux2_1_A0 hold313/A m_blake2.m_hash256.h_flat\[192\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout374/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold353/X fanout580/X
+ VGND VGND VPWR VPWR hold354/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1/Y
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ sky130_fd_sc_hd__nand2b_2
Xm_blake2.m_hash256.m_matrix\[9\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold585/X hold750/A fanout575/X VGND VGND VPWR VPWR hold586/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[20\]_sky130_fd_sc_hd__mux2_1_A1_S fanout218/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__inv_2_Y
+ fanout478/X VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/A
+ sky130_fd_sc_hd__inv_2
Xm_blake2.m_hash256.m_matrix\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold551/X fanout546/X
+ VGND VGND VPWR VPWR hold552/A sky130_fd_sc_hd__mux2_1
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_1278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[3\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1153/X hold1198/A fanout582/X VGND VGND VPWR VPWR hold1154/A sky130_fd_sc_hd__mux2_1
XFILLER_29_1174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold345/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_18_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1001/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[10\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__xnor2_2_A hold1089/A hold377/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[3\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold279/X fanout409/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X/B2 m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X/B2
+ fanout557/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.h_flat\[196\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold103/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_52_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1239/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold541/A fanout145/X fanout97/X m_blake2.m_hash256.m_matrix\[6\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout244_A fanout248/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_43_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[10\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B/C
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.v_q\[2\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold452/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout509_A fanout539/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__or2_2_A hold238/A fanout248/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout411_A fanout412/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[1\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_B
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_fanout499_X fanout499/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xdata\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X m_io.m_config.data_i\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ hold9/X fanout308/X VGND VGND VPWR VPWR data\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[25\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__a22o_2_A1 hold599/A fanout293/X
+ fanout286/X hold709/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold906/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold731/X m_blake2.m_hash256.v_q\[15\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout209/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_43_1116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1234/X fanout228/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold248/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0 hold458/A m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout389/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_1436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold1042/X fanout164/X m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__or2_2_A/X fanout617/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[35\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_16_737 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B/X
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2b_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X
+ hold1067/A fanout130/X fanout122/X m_blake2.m_hash256.m_matrix\[15\]\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_31_729 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1114/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__and2_2_B fanout435/X hold600/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_15_1207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload16/A m_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.h_flat\[119\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0
+ m_blake2.m_hash256.h_flat\[170\]_sky130_fd_sc_hd__and3_2_C/X m_blake2.m_hash256.v_q\[5\]\[2\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/Y
+ fanout513/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[162\]_sky130_fd_sc_hd__a21o_2_A1/B1
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold774/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__mux2_1_A0 hold506/X m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout414/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[17\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XFILLER_79_921 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[3\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout258/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[205\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold64/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__xor2_2_A hold1044/A hold287/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[17\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_A m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[23\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A1
+ fanout239/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[214\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold191/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.d_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_1165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[15\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1201/X m_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout565/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_692 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__mux2_1_A0 hold283/X m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout229/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_47_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkload24/A m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold473/A sky130_fd_sc_hd__dfxtp_1
XFILLER_37_1443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__xor2_2_B hold628/A hold403/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout349/X m_blake2.m_hash256.v_q\[5\]\[8\]_sky130_fd_sc_hd__a22o_2_A1/X fanout178/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
Xhold903 hold903/A VGND VGND VPWR VPWR hold903/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold914 hold914/A VGND VGND VPWR VPWR hold914/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold936 hold936/A VGND VGND VPWR VPWR hold936/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 hold925/A VGND VGND VPWR VPWR hold925/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[11\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.v_q\[11\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1182/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold347/A m_blake2.m_hash256.h_flat\[218\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout369/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold958 hold958/A VGND VGND VPWR VPWR hold958/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 hold947/A VGND VGND VPWR VPWR hold947/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold969 hold969/A VGND VGND VPWR VPWR hold969/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkload29_A clkload29/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout63/X fanout75/X
+ hold1253/A m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[3\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold411/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A fanout194/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A0 hold329/A m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout532/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1001/A fanout26/X fanout54/X hold1167/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout361_A fanout361/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A_A m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_873 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A/C
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1/Y
+ sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout195/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1170/A fanout82/X fanout70/X hold1200/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_52_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.d_q\[23\]_sky130_fd_sc_hd__xor2_2_A_B m_blake2.m_hash256.m_g.a_q\[23\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_386 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_718 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[1\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_19_clk/X
+ m_blake2.m_hash256.m_matrix\[1\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1088/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload34/A m_blake2.m_hash256.v_q\[5\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold548/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout183/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_2
XANTENNA_fanout414_X fanout414/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__and2_2_A_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_751 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__mux2_1_A0 hold628/X m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout234/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[2\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_75_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold623/X m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout160/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_699 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X m_blake2.m_hash256.h_flat\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold83/A sky130_fd_sc_hd__dfxtp_1
XFILLER_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1
+ m_io.m_config.data_i\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold788/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_48_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__xnor2_2_A hold670/A hold813/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[1\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkload22/A m_blake2.m_hash256.m_g.a0\[22\]_sky130_fd_sc_hd__xor2_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_44_832 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_44_810 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_884 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__mux2_1_A0/X
+ m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__or2_2_B/B fanout318/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.h_flat\[24\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XFILLER_71_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold1069/X fanout203/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold403/X m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout414/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout94/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_887 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1 m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B
+ fanout358/X fanout262/X m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__and3_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[5\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_54_1020 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_773 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout155/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_1097 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2/X m_blake2.m_hash256.v_q\[0\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__and2_2_A/B sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold968/A fanout24/X fanout40/X hold515/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_8_744 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_755 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__and2_2_B fanout441/X hold264/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[180\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_16_clk/X
+ hold639/X VGND VGND VPWR VPWR hold638/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/B1_N
+ m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1/A2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nor2_2
XFILLER_32_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[11\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold845/X hold1175/A fanout552/X VGND VGND VPWR VPWR hold846/A sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold262/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_B
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A m_blake2.m_hash256.g_buffer\[23\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[23\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A0 hold119/A m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_72_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[16\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout22/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__or2_2_A hold1228/A fanout388/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_26_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A0 hold116/A m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_1035 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout229/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__or2_2_A hold1114/A fanout394/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[29\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XFILLER_39_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_1188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.h_flat\[50\]_sky130_fd_sc_hd__nor2_2_B_A fanout484/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1 m_blake2.m_hash256.m_g.d_q\[30\]_sky130_fd_sc_hd__xor2_2_A/B
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/B m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ sky130_fd_sc_hd__a21oi_1
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[7\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold821/A sky130_fd_sc_hd__dfxtp_1
XFILLER_35_821 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold200/A m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout530/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold802/X m_blake2.m_hash256.g_y_buf\[27\]_sky130_fd_sc_hd__o32a_2_X/B2 fanout578/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_74_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_37_clk/X m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[4\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_50_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_802 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold515/A fanout88/X fanout144/X hold629/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_37_1273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2/X
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a2111o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__o211a_2
XTAP_TAPCELL_ROW_79_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__or2_2_B fanout498/X hold57/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[207\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B_A fanout437/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout207_A fanout208/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y
+ m_blake2.m_hash256.m_g.b_q\[24\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold711 hold711/A VGND VGND VPWR VPWR hold711/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N
+ m_blake2.m_hash256.m_matrix\[0\]\[7\]_sky130_fd_sc_hd__o22ai_2_A1/Y m_blake2.m_hash256.v_q\[0\]\[7\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3_2_B/A
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__dfxtp_2_Q clkload11/A m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold138/A sky130_fd_sc_hd__dfxtp_1
Xhold700 hold700/A VGND VGND VPWR VPWR hold700/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold755 hold755/A VGND VGND VPWR VPWR hold755/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold733 hold733/A VGND VGND VPWR VPWR hold733/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_38_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold722 hold722/A VGND VGND VPWR VPWR hold722/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 hold744/A VGND VGND VPWR VPWR hold744/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[9\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1196/A sky130_fd_sc_hd__dfxtp_1
Xhold788 hold788/A VGND VGND VPWR VPWR hold788/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 hold777/A VGND VGND VPWR VPWR hold777/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 hold766/A VGND VGND VPWR VPWR hold766/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[7\]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1
+ fanout269/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold1228/X m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout156/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold799 hold799/A VGND VGND VPWR VPWR hold799/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_33_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__a311o_2_A1 hold1129/A fanout355/X
+ fanout249/X m_blake2.m_hash256.v_q\[11\]\[19\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.v_q\[10\]\[19\]_sky130_fd_sc_hd__o21a_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[19\]_sky130_fd_sc_hd__o22a_2_X/B1
+ sky130_fd_sc_hd__a311o_1
XFILLER_69_250 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout197_X fanout197/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_935 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_buffer\[8\].m_c_buf m_blake2.m_hash256.g_buffer\[8\].m_c_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[8\].m_c_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_57_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_1108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__a211oi_2_A1 hold562/A fanout281/X
+ m_blake2.m_hash256.v_q\[1\]\[31\]_sky130_fd_sc_hd__a22o_2_A1/X fanout390/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[31\]_sky130_fd_sc_hd__a211oi_2_A1/Y
+ sky130_fd_sc_hd__a211oi_1
Xm_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__a31o_2_A3 fanout472/X fanout476/X
+ hold340/A fanout363/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A_B
+ m_blake2.m_hash256.block_idx_plus_one_q\[46\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_48_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_824 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_40_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_A1
+ fanout290/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__a31o_2_A3 fanout447/X fanout480/A
+ hold142/A fanout532/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[236\]_sky130_fd_sc_hd__a31o_2_A3/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_m_io.m_config.ll_q\[40\]_sky130_fd_sc_hd__and3_2_A_B fanout465/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[0\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[5\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold778/X m_blake2.m_hash256.m_matrix\[6\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout553/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A0 ANTENNA_5/DIODE m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout501/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[8\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload15/A m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.data_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.block_idx_plus_one_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.block_idx_plus_one_q\[7\]_sky130_fd_sc_hd__and4_2_C/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
Xm_blake2.m_hash256.m_matrix\[6\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[6\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold346/A sky130_fd_sc_hd__dfxtp_1
Xhold82 hold82/A VGND VGND VPWR VPWR hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.d_q\[31\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
Xhold71 hold71/A VGND VGND VPWR VPWR hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B
+ fanout401/X m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold93 hold93/A VGND VGND VPWR VPWR hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout413/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[53\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1
+ fanout421/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y
+ fanout228/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout290/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold1005/A fanout135/X fanout118/X hold1169/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.c_q\[31\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_14_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold1086/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[1\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout126/X fanout150/X
+ hold706/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[8\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A hold559/X
+ VGND VGND VPWR VPWR hold558/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__and3_2_A hold614/A fanout465/X fanout373/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[51\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XFILLER_32_1170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 ANTENNA_2/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X hold529/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o41a_2_B1
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1/Y
+ m_blake2.m_hash256.m_g.b_q\[8\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B/X
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__o41a_1
Xm_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[219\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xfanout509 fanout539/X VGND VGND VPWR VPWR fanout509/X sky130_fd_sc_hd__buf_2
XFILLER_80_1422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[23\]_sky130_fd_sc_hd__a211o_2_A1_A2 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold247/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[136\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[20\]_sky130_fd_sc_hd__a221o_2_B2_B1 fanout307/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_651 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A hold337/A m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout178/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_1237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout157_A fanout160/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1000/X fanout568/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xor2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__and2_2_B fanout433/X hold202/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[139\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[13\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout31/X fanout39/X
+ hold974/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2
+ m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__mux2_1_A1/X m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ fanout511/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ sky130_fd_sc_hd__a21bo_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout290/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[8\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0
+ m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__xnor2_2_A hold432/A hold1207/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout112_X fanout112/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold530 hold530/A VGND VGND VPWR VPWR hold530/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_A1
+ fanout286/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[28\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold563 hold563/A VGND VGND VPWR VPWR hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 hold552/A VGND VGND VPWR VPWR hold552/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold541 hold541/A VGND VGND VPWR VPWR hold541/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold585 hold585/A VGND VGND VPWR VPWR hold585/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 hold596/A VGND VGND VPWR VPWR hold596/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold574 hold574/A VGND VGND VPWR VPWR hold574/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_A
+ m_io.m_config.kk_q\[5\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_A2
+ m_blake2.m_hash256.m_g.b_q\[13\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__xnor2_2_B hold742/A hold441/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[13\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold1241 hold1241/A VGND VGND VPWR VPWR hold1241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1252 hold1252/A VGND VGND VPWR VPWR hold1252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1230 hold1230/A VGND VGND VPWR VPWR hold1230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1263 hold1263/A VGND VGND VPWR VPWR hold1263/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__xnor2_2_A hold567/A hold512/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[18\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__xnor2_2_B_A
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2/A1_N
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_813 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__nand2b_2_B_B m_blake2.m_hash256.m_g.m_add_1.x2_i\[8\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__or2_2_A m_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__or2_2_A/A
+ fanout241/X VGND VGND VPWR VPWR m_io.m_config.ll_q\[1\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X
+ hold1183/A fanout114/X m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ fanout106/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A1
+ sky130_fd_sc_hd__a2111o_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout294/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.kk_q\[3\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload26/A m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[13\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__or2_2_B_A fanout485/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.res_cnt_q\[4\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/B sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_A0 m_blake2.m_hash256.v_q\[15\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1 m_blake2.m_hash256.g_y_buf\[5\]_sky130_fd_sc_hd__o22a_2_X/A1
+ fanout100/X m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/B1
+ m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/B2 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1/Y sky130_fd_sc_hd__o22ai_4
Xclkbuf_3_3_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkload1/A sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_44_clk/X
+ m_blake2.m_hash256.h_flat\[143\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold30/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[11\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout574/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[11\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_buffer\[9\].m_y_buf m_blake2.m_hash256.g_buffer\[9\].m_y_buf/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[9\].m_y_buf/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_C1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__xnor2_2_A hold1129/A hold557/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_5_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__a31o_2_B1_B1
+ m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[152\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold632/X fanout327/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[144\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[13\]\[27\]_sky130_fd_sc_hd__nor2_2_A hold1024/A fanout375/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__a221o_2_B2/C1 sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold558/X fanout572/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_1300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.res_cnt_q\[2\]_sky130_fd_sc_hd__nor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout157/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[8\]_sky130_fd_sc_hd__xor2_2_X/A sky130_fd_sc_hd__nand2_1
XFILLER_1_794 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/B
+ sky130_fd_sc_hd__xor2_4
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_S fanout303/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A
+ m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y/A m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_49_787 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_1090 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B fanout495/X hold146/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[78\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[15\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/A
+ m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
XFILLER_17_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.ll_q\[59\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__a221o_2_B2_C1 fanout269/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_665 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__xnor2_2_A hold301/A hold965/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ hold303/A fanout306/X m_blake2.m_hash256.v_q\[12\]\[29\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[29\]_sky130_fd_sc_hd__nor2_2_Y/B sky130_fd_sc_hd__a21oi_1
XFILLER_34_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xor2_2
Xm_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[26\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ sky130_fd_sc_hd__a21o_1
XFILLER_30_1129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[3\]_sky130_fd_sc_hd__and3_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[222\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A0 hold412/A m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout520/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
Xfanout339 fanout340/X VGND VGND VPWR VPWR fanout339/X sky130_fd_sc_hd__clkbuf_4
Xfanout328 fanout330/X VGND VGND VPWR VPWR fanout328/X sky130_fd_sc_hd__buf_4
Xfanout317 fanout342/A VGND VGND VPWR VPWR fanout317/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1140/A fanout126/X fanout142/X hold865/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xfanout306 fanout307/X VGND VGND VPWR VPWR fanout306/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__or2_2_A hold305/A fanout378/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[28\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_52_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_A1
+ fanout255/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__xnor2_2_A hold296/A m_blake2.m_hash256.v_q\[14\]\[21\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout274_A fanout274/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_713 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_54_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[46\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_65_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1053/A fanout116/X fanout121/X m_blake2.m_hash256.m_matrix\[15\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[22\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[4\]_sky130_fd_sc_hd__xor2_2_X/X
+ sky130_fd_sc_hd__xor2_1
XFILLER_74_1012 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X
+ m_blake2.m_hash256.h_flat\[169\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold102/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_fanout441_A fanout442/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout327_X fanout327/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__mux2_1_A1_S fanout215/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_8_clk/X m_blake2.m_hash256.h_flat\[82\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X
+ m_blake2.m_hash256.v_q\[7\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold805/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X
+ m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__mux2_1_A0 hold349/A hash\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ fanout392/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold360 hold360/A VGND VGND VPWR VPWR hold360/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 hold371/A VGND VGND VPWR VPWR hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[91\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold155/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[83\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold393 hold393/A VGND VGND VPWR VPWR hold393/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 hold382/A VGND VGND VPWR VPWR hold382/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_d\[28\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2
+ m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A hash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_5_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_S fanout415/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold752/X fanout585/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[15\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xnor2_2_A_A
+ m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/X VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xhold1060 hold1060/A VGND VGND VPWR VPWR hold1060/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[20\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhash\[2\]_sky130_fd_sc_hd__mux2_1_A1 hash\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0 hash\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout430/X VGND VGND VPWR VPWR hash\[2\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
Xhold1082 hold1082/A VGND VGND VPWR VPWR hold1082/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_46_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1093 hold1093/A VGND VGND VPWR VPWR hold1093/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1071 hold1071/A VGND VGND VPWR VPWR hold1071/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_25_clk/X
+ m_blake2.m_hash256.v_q\[13\]\[9\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold1218/A sky130_fd_sc_hd__dfxtp_1
XFILLER_61_727 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B fanout496/X hold187/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[43\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[24\]_sky130_fd_sc_hd__a22o_2_A1_A2 fanout190/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1156/X m_blake2.m_hash256.m_matrix\[12\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout550/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__xor2_2_X
+ fanout467/X fanout475/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__xor2_4
Xm_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A0 hold128/A m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout514/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_A_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y/C
+ m_blake2.m_hash256.m_g.a0\[19\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X/A
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_13_clk/X
+ m_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[14\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A hold673/A m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[7\]_sky130_fd_sc_hd__xor2_2_A/X
+ sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout110/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[8\]_sky130_fd_sc_hd__a211oi_2_A1_A2 fanout284/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0 m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A/Y
+ hold68/A fanout428/X VGND VGND VPWR VPWR m_io.m_config.kk_q\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1112/X
+ fanout565/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_1236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[27\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[28\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C/Y
+ sky130_fd_sc_hd__nand3_1
XFILLER_29_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_Y m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkload13/A m_blake2.m_hash256.m_matrix\[9\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold696/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_hash\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1 hash\[6\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout62/X fanout42/X
+ hold1058/A m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[8\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout181/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold729/A fanout134/X fanout143/X hold757/A m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XFILLER_32_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[13\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout44/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[18\]_sky130_fd_sc_hd__mux2_1_A0_S fanout212/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D/A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C/Y
+ VGND VGND VPWR VPWR fanout127/A sky130_fd_sc_hd__and4_2
XTAP_TAPCELL_ROW_41_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold629/A fanout52/X fanout68/X hold1208/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_1371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_54_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout103 fanout103/A VGND VGND VPWR VPWR fanout103/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand3_2_C
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1/A2
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand3_2_C/B
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[16\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1/A2
+ sky130_fd_sc_hd__nand3_1
XANTENNA_fanout489_A fanout500/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout147 fanout147/A VGND VGND VPWR VPWR fanout147/X sky130_fd_sc_hd__clkbuf_2
Xfanout136 fanout139/X VGND VGND VPWR VPWR fanout136/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout391_A fanout398/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout114 fanout115/A VGND VGND VPWR VPWR fanout114/X sky130_fd_sc_hd__clkbuf_4
Xfanout125 fanout127/A VGND VGND VPWR VPWR fanout125/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_860 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout158 fanout160/A VGND VGND VPWR VPWR fanout158/X sky130_fd_sc_hd__buf_2
XFILLER_41_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout169 fanout170/A VGND VGND VPWR VPWR fanout169/X sky130_fd_sc_hd__buf_4
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_S fanout419/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1093 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_47_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A1
+ m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[5\]_sky130_fd_sc_hd__xnor2_2_Y/B
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_io.m_config.ll_q\[58\]_sky130_fd_sc_hd__and3_2_A_B fanout463/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_757 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1118 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_76_1107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[18\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout181/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_1099 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_919 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_48_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_A
+ fanout408/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[8\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1131/X m_blake2.m_hash256.m_matrix\[8\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout593/X
+ VGND VGND VPWR VPWR hold1132/A sky130_fd_sc_hd__mux2_1
XFILLER_54_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout148/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A/X
+ m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[6\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ sky130_fd_sc_hd__nand2b_2
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X/A1
+ m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X/A2 m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X/B1
+ fanout181/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout92_X fanout92/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ sky130_fd_sc_hd__a21o_1
Xhold190 hold190/A VGND VGND VPWR VPWR hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[14\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout64/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_893 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nor2_2_Y
+ fanout466/X fanout469/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X/B
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_53_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold557/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[4\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_1117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold629/X fanout552/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[20\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_771 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_955 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[11\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[11\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold503/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[12\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X
+ m_blake2.m_hash256.v_q\[12\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold907/A sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_690 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout150/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_1268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_661 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[12\]\[1\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1194/X fanout225/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[12\]\[1\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X
+ m_blake2.m_hash256.m_g.c_q\[16\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[17\]_sky130_fd_sc_hd__nand3_2_A/B
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X/A
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X/B
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/B
+ sky130_fd_sc_hd__or3_4
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_26_clk/X
+ m_blake2.m_hash256.v_q\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold419/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout231/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_1039 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold1098/X m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout298/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[13\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_863 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout91/X
+ fanout119/X hold1197/A m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_37_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__or2_2_A hold731/A fanout369/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[10\]_sky130_fd_sc_hd__or2_2_A/X
+ sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__mux2_1_A0 hold644/X m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout300/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A/Y
+ m_blake2.m_hash256.v_q\[11\]\[2\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[7\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/A0 sky130_fd_sc_hd__xnor2_2
XFILLER_80_888 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_782 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_1195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout237_A fanout239/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_977 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout86/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_31_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout404_A fanout406/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21bo_2_X
+ hold1180/X fanout152/X fanout482/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a21bo_1
Xm_blake2.m_hash256.m_matrix\[15\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[15\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold840/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1
+ fanout194/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[30\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout176/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1231/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout192/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout200/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[26\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_A
+ fanout401/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0 hold468/X m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[22\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold358/A sky130_fd_sc_hd__dfxtp_1
XFILLER_58_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N_Y m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__nand3b_2_A_N/Y
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[3\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold458/X fanout411/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[7\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold820/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o31a_2_A3
+ fanout453/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or3_2_A_1/X
+ m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A/B
+ sky130_fd_sc_hd__o31a_1
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1
+ fanout181/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold342/X m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout160/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_70_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_1322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[4\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold900/X hold890/X fanout553/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[4\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold466/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X
+ m_io.m_block_data.data_cnt_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold2/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__o21a_2_A1 m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B/A
+ fanout364/X fanout169/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[18\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N
+ m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N/X
+ sky130_fd_sc_hd__and2b_1
Xm_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[187\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[195\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1
+ fanout468/X fanout401/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/X
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1/X m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1/X
+ sky130_fd_sc_hd__a311o_1
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1 m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR fanout239/A sky130_fd_sc_hd__or2_2
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[22\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[2\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[22\]_sky130_fd_sc_hd__or2_2_A/B sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1 m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A/A
+ fanout459/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A/C fanout444/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_1/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout419/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_1331 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__or2_2_A hold461/A fanout245/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[15\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[10\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout54/X
+ fanout78/X m_blake2.m_hash256.m_matrix\[8\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[14\]_sky130_fd_sc_hd__mux2_1_A0_S fanout155/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__mux2_1_A0_S fanout157/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold382/A m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout517/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B/Y m_blake2.m_hash256.v_q\[2\]\[16\]_sky130_fd_sc_hd__xor2_2_B/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[0\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ hold484/X VGND VGND VPWR VPWR hold483/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.v_q\[4\]\[24\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold703/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[28\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout68/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[18\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_4
XFILLER_24_1050 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__mux2_1_A0 hold68/A m_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout503/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[9\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_37_1466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_752 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[2\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_12_clk/X
+ m_blake2.m_hash256.m_matrix\[2\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold970/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkload18/A m_blake2.m_hash256.v_q\[6\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold396/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__mux2_1_A0 hold479/X m_blake2.m_hash256.v_q\[3\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_970 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold904 hold904/A VGND VGND VPWR VPWR hold904/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_77_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold926 hold926/A VGND VGND VPWR VPWR hold926/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 hold915/A VGND VGND VPWR VPWR hold915/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 hold937/A VGND VGND VPWR VPWR hold937/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold347/X fanout213/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold948 hold948/A VGND VGND VPWR VPWR hold948/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ hold594/X fanout201/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xhold959 hold959/A VGND VGND VPWR VPWR hold959/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__and3_2_A hold240/A fanout464/X fanout383/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__and3_2_A/X sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_36_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.h_flat\[211\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold451/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold969/X fanout568/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1
+ fanout284/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[0\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.h_flat\[48\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2
+ fanout289/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_d\[3\]_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__o21a_2_X_B1
+ fanout185/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A fanout189/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2
+ fanout290/X m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[72\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2/Y
+ sky130_fd_sc_hd__a21boi_1
Xm_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[220\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold329/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[212\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__a22o_2_A1 hold123/X fanout327/X
+ m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__a22o_2_A1/B1 fanout520/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[248\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2
+ fanout404/X m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.v_q\[2\]\[6\]_sky130_fd_sc_hd__a211o_2_A1/X
+ m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2/A2_N
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__mux2_1_A0 hold284/X m_blake2.m_hash256.v_q\[7\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ fanout232/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[31\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[8\]\[26\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold941/A sky130_fd_sc_hd__dfxtp_1
XFILLER_38_885 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[4\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_4_clk/X
+ m_blake2.m_hash256.m_matrix\[4\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold900/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__a31o_2_A3_A1 fanout472/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout354_A fanout361/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkload29/A m_blake2.m_hash256.v_q\[4\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold393/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_2
XFILLER_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold998/X fanout586/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout521_A fanout524/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout142_X fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[8\]\[27\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1191/X fanout224/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[27\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_741 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__and2_2_A_B m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_hash\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S fanout314/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_763 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__and2_2_A/B
+ fanout424/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_7_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_785 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout407_X fanout407/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B1
+ m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[4\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold883/X hold1078/A fanout547/X VGND VGND VPWR VPWR hold884/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[4\]_sky130_fd_sc_hd__mux2_1_A0_S fanout236/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[10\]\[1\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold281/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_0_clk/X
+ m_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[6\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.g_b\[5\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2_A1 m_io.m_config.ll_q\[34\]_sky130_fd_sc_hd__a22oi_2_B2/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y/Y VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[26\]_sky130_fd_sc_hd__xor2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X
+ fanout258/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.round_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_23_clk/X m_blake2.m_hash256.round_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout458/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold693/X fanout556/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__o21a_2_A1 hold979/A fanout387/X
+ fanout172/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[22\]_sky130_fd_sc_hd__o21a_2_A1/X
+ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_8_Left_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout128/X fanout96/X
+ m_blake2.m_hash256.m_matrix\[6\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout196/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout188/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[25\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2/X
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A/B
+ sky130_fd_sc_hd__or2_1
XFILLER_5_1442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/A sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or2_2_B
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A/C
+ sky130_fd_sc_hd__or2_1
XFILLER_44_844 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold631/X fanout573/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[19\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_71_696 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold924/A fanout58/X fanout38/X hold690/A m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[24\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_34_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload12/A m_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold662/X fanout566/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[7\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_1330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[6\]_sky130_fd_sc_hd__and2b_2_B_A_N m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N/A
+ m_blake2.m_hash256.m_g.a_q\[5\]_sky130_fd_sc_hd__and3_2_A/X m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N/X
+ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_22_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_40_clk/X
+ m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold58/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__or2_2_B_A fanout499/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X
+ hold486/A fanout100/X m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B1
+ m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ sky130_fd_sc_hd__o22a_2
Xm_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_61_clk/X
+ m_blake2.m_hash256.h_flat\[116\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold126/A sky130_fd_sc_hd__dfxtp_1
Xdata_idx\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X hold4/X VGND VGND VPWR
+ VPWR data_idx\[3\]_sky130_fd_sc_hd__and4_2_A/B sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.g_b\[14\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_72_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold119/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.v_q\[0\]\[0\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_72_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__nand2_2_B fanout439/X hold278/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[229\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
Xm_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ hold876/A fanout118/X fanout94/X hold1031/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[125\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold116/X fanout324/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[117\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_79_785 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B_A
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_1156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold585/A fanout33/X fanout40/X m_blake2.m_hash256.m_matrix\[14\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[23\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_446 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_38_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[3\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload8/A m_blake2.m_hash256.m_matrix\[3\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold400/A sky130_fd_sc_hd__dfxtp_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D_sky130_fd_sc_hd__a22o_2_X m_io.m_config.data_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ m_io.cmd\[4\]_sky130_fd_sc_hd__and2b_2_B/X uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1
+ hash\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A1_S fanout409/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[194\]_sky130_fd_sc_hd__and2_2_B_A fanout430/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1/X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2/Y
+ sky130_fd_sc_hd__o21ai_4
Xm_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[38\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold200/X fanout332/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold627/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[30\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_73_clk clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_73_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[20\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_6_clk/X
+ m_blake2.m_hash256.m_matrix\[5\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1177/A sky130_fd_sc_hd__dfxtp_1
XFILLER_34_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__and3_2_B/X m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[56\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XFILLER_61_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and3_2_C
+ m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B/A fanout445/X
+ m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X/B VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__o21a_2_A1/A2
+ sky130_fd_sc_hd__and3_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[6\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1
+ fanout404/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_1187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold246/X fanout163/X m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__or2_2_A/X fanout613/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XFILLER_30_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_20_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__and2_2_B fanout433/X hold66/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[240\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold1037/A sky130_fd_sc_hd__dfxtp_1
Xuo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X hash\[0\]_sky130_fd_sc_hd__or2_2_B/B
+ uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X/B1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X/B1
+ VGND VGND VPWR VPWR uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7/D sky130_fd_sc_hd__a21o_1
Xhold712 hold712/A VGND VGND VPWR VPWR hold712/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B fanout438/X hold93/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[107\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xhold701 hold701/A VGND VGND VPWR VPWR hold701/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A0 hold265/A m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout532/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout102_A fanout103/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold723 hold723/A VGND VGND VPWR VPWR hold723/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold734 hold734/A VGND VGND VPWR VPWR hold734/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 hold745/A VGND VGND VPWR VPWR hold745/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_io.m_config.ll_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1240/A sky130_fd_sc_hd__dfxtp_1
Xhold756 hold756/A VGND VGND VPWR VPWR hold756/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 hold778/A VGND VGND VPWR VPWR hold778/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold767 hold767/A VGND VGND VPWR VPWR hold767/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__o21a_2_A1 m_blake2.m_hash256.v_q\[9\]\[15\]_sky130_fd_sc_hd__xor2_2_A/A
+ fanout386/X fanout251/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[15\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A0 hold56/A m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout528/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xhold789 hold789/A VGND VGND VPWR VPWR hold789/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_925 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__o21a_2_A1_B1 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.block_idx_plus_one_q\[24\]_sky130_fd_sc_hd__and3_2_B/C m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__o21ai_2_A1/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout471_A fanout472/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B fanout429/X hold38/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[40\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__xnor2_2_A hold279/A m_blake2.m_hash256.v_q\[8\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_811 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q_Q
+ m_blake2.m_hash256.v_q\[13\]\[1\]_sky130_fd_sc_hd__a221o_2_A1/B2 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_64_clk clkload2/A VGND VGND VPWR VPWR clkload24/A sky130_fd_sc_hd__clkbuf_8
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout524_X fanout524/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_836 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B/A
+ m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[21\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/A
+ sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X
+ fanout299/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
Xm_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/B VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X/X
+ sky130_fd_sc_hd__xor2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1
+ fanout252/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_1358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2
+ fanout172/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[200\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[208\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[1\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[9\]\[21\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[14\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[55\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X
+ hold930/A fanout98/X fanout122/X hold948/A m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[2\]_sky130_fd_sc_hd__o32a_2_B2/A2
+ sky130_fd_sc_hd__a221o_1
XFILLER_49_1145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_1301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[64\]_sky130_fd_sc_hd__mux2_1_A0/X
+ ANTENNA_5/DIODE fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[56\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_1465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_B2
+ fanout288/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[77\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1
+ fanout283/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C block_last_sky130_fd_sc_hd__a32o_2_B2/A3
+ m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B hold652/A VGND VGND VPWR
+ VPWR m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/Y sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__nor2_2_B fanout499/X hold1022/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[246\]_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
Xhold72 hold72/A VGND VGND VPWR VPWR hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A VGND VGND VPWR VPWR hold83/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold94 hold94/A VGND VGND VPWR VPWR hold94/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__xnor2_2_A hold251/A hold714/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[19\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_3_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold1188/A fanout124/X fanout120/X hold648/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_55_clk clkload3/A VGND VGND VPWR VPWR clkload28/A sky130_fd_sc_hd__clkbuf_8
XTAP_TAPCELL_ROW_80_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X
+ hold350/A fanout351/X fanout183/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_27_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1053/X
+ fanout563/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_66_clk/X
+ m_blake2.m_hash256.v_q\[2\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold524/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_30_clk/X m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold642/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_14_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A0 hold90/A m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout535/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y
+ fanout47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[26\]_sky130_fd_sc_hd__inv_2_Y/Y sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_74_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_3 ANTENNA_3/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__a32o_2_A1_A2 fanout346/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold563/A fanout59/X fanout75/X hold863/A m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XANTENNA_m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y
+ m_blake2.m_hash256.g_b\[23\]_sky130_fd_sc_hd__inv_2_Y/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.c_q\[19\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout96/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A0 hold50/A m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout526/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B
+ fanout477/X m_blake2.m_hash256.v_q\[10\]\[30\]_sky130_fd_sc_hd__and3_2_B/C VGND
+ VGND VPWR VPWR fanout254/A sky130_fd_sc_hd__nor2_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[23\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_A2
+ m_blake2.m_hash256.v_q\[15\]\[23\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload30/A
+ m_blake2.m_hash256.block_idx_plus_one_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR hold1245/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout127/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__xnor2_2_B hold1166/A hold740/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[16\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold498/X m_blake2.m_hash256.m_g.d_q\[22\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ fanout419/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[3\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_hash\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_Q hash\[7\]_sky130_fd_sc_hd__and2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y
+ fanout238/X m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[12\]_sky130_fd_sc_hd__a21oi_2_Y/B1 sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_46_clk clkload5/A VGND VGND VPWR VPWR clkload34/A sky130_fd_sc_hd__clkbuf_8
XFILLER_62_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_35_663 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_803 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold876/A fanout30/X fanout38/X hold794/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[16\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_g.d_q\[18\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A/B
+ hold655/X fanout410/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_34_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_847 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1060 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B
+ m_blake2.m_hash256.v_q\[11\]\[8\]_sky130_fd_sc_hd__mux2_1_A1/A0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y
+ fanout237/X m_blake2.m_hash256.v_q\[13\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/X m_blake2.m_hash256.v_q\[15\]\[26\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[26\]_sky130_fd_sc_hd__nor2_2_Y/A sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[15\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout63/X
+ fanout71/X m_blake2.m_hash256.m_matrix\[7\]\[18\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND
+ VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[18\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/B1
+ sky130_fd_sc_hd__a22o_1
XFILLER_31_891 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout317_A fanout342/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold520 hold520/A VGND VGND VPWR VPWR hold520/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold531 hold531/A VGND VGND VPWR VPWR hold531/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold553 hold553/A VGND VGND VPWR VPWR hold553/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or3_2_A
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[25\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.m_g.c_q\[27\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or3_2_A/X
+ sky130_fd_sc_hd__or3_1
Xm_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__xor2_2_B hold776/A hold735/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[8\]_sky130_fd_sc_hd__xor2_2_B/X sky130_fd_sc_hd__xor2_1
Xhold542 hold542/A VGND VGND VPWR VPWR hold542/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_57_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout34/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold586 hold586/A VGND VGND VPWR VPWR hold586/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 hold597/A VGND VGND VPWR VPWR hold597/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 hold564/A VGND VGND VPWR VPWR hold564/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 hold575/A VGND VGND VPWR VPWR hold575/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/A1
+ m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/A2 m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/B1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[11\]_sky130_fd_sc_hd__a21oi_2_Y/Y sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[0\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout18/X hold134/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[0\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
Xm_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ m_blake2.m_hash256.m_matrix\[7\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout108/X fanout121/X
+ hold867/A m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[6\]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
XFILLER_58_711 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold1220 hold1220/A VGND VGND VPWR VPWR hold1220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1231 hold1231/A VGND VGND VPWR VPWR hold1231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1242 hold1242/A VGND VGND VPWR VPWR hold1242/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_A_sky130_fd_sc_hd__o21a_2_X
+ m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or3_2_A_2/C m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__or3_2_A/C
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o41a_2_A2/B1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D/A
+ sky130_fd_sc_hd__o21a_1
Xhold1253 hold1253/A VGND VGND VPWR VPWR hold1253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1264 hold1264/A VGND VGND VPWR VPWR hold1264/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_37_clk clkload5/A VGND VGND VPWR VPWR clkbuf_leaf_37_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_2
XFILLER_22_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A
+ m_blake2.m_hash256.g_buffer\[26\].m_y_buf/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X/A
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A/B
+ sky130_fd_sc_hd__xor2_1
Xm_blake2.m_hash256.v_q\[14\]\[5\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__xnor2_2_A/B
+ m_blake2.m_hash256.v_q\[15\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout210/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_24_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout18_X fanout18/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout293/X m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[99\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2/X
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_matrix\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_3_clk/X
+ m_blake2.m_hash256.m_matrix\[3\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1003/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A0 hold1102/A m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout505/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_33_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[36\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y
+ hold317/X fanout304/X m_blake2.m_hash256.v_q\[12\]\[10\]_sky130_fd_sc_hd__a221o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[10\]_sky130_fd_sc_hd__nor2_2_Y/B sky130_fd_sc_hd__a21oi_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[1\]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout82/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_S fanout155/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y fanout342/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__dfxtp_2_Q_Q fanout465/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_1429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[6\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout286/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y
+ hold308/A fanout375/X fanout185/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[27\]_sky130_fd_sc_hd__a21oi_2_Y/A1
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21o_2_A1
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[18\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1/X
+ m_blake2.m_hash256.m_g.d_q\[3\]_sky130_fd_sc_hd__xor2_2_A/X VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/B
+ sky130_fd_sc_hd__a21o_1
XFILLER_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[26\]_sky130_fd_sc_hd__a32o_2_A1_B1 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1/Y m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[30\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_2
Xm_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__xnor2_2_A hold1069/A hold485/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[24\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_28_clk clkload1/A VGND VGND VPWR VPWR clkbuf_leaf_28_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.m_g.d_q\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload29/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__xnor2_2_A m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__inv_2_A/A
+ m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR m_io.m_config.nn_q\[2\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B
+ m_io.m_config.cfg_cnt_q\[1\]_sky130_fd_sc_hd__or3_2_A/X m_io.m_config.nn_q\[0\]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor2_2_Y/B
+ VGND VGND VPWR VPWR m_io.m_config.nn_q\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X/A2
+ sky130_fd_sc_hd__or2_2
XFILLER_60_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_685 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[33\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N
+ m_blake2.m_hash256.block_idx_plus_one_q\[34\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__nor2_2_B
+ fanout367/X m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[2\]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_32_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.v_q\[13\]\[10\]_sky130_fd_sc_hd__a221o_2_A1_B1 fanout260/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_873 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_895 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_47_clk_A clkload4/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[158\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold412/X fanout328/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[150\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_1015 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout329 fanout330/X VGND VGND VPWR VPWR fanout329/X sky130_fd_sc_hd__buf_2
Xfanout307 fanout307/A VGND VGND VPWR VPWR fanout307/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y/B
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y/B
+ sky130_fd_sc_hd__nand3_1
Xm_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a31o_2_X
+ m_blake2.m_hash256.g_b\[8\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B/Y
+ m_blake2.m_hash256.m_g.a0\[10\]_sky130_fd_sc_hd__xnor2_2_Y/A m_blake2.m_hash256.m_g.a0\[9\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A/X
+ m_blake2.m_hash256.g_b\[9\]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[11\]_sky130_fd_sc_hd__xnor2_2_Y/A
+ sky130_fd_sc_hd__a31o_1
Xfanout318 fanout323/X VGND VGND VPWR VPWR fanout318/X sky130_fd_sc_hd__clkbuf_4
Xm_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1 fanout446/X fanout478/X
+ fanout507/X VGND VGND VPWR VPWR fanout342/A sky130_fd_sc_hd__a21oi_4
XTAP_TAPCELL_ROW_52_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[29\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout286/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_725 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_19_clk clkbuf_3_2_0_clk/X VGND VGND VPWR VPWR clkbuf_leaf_19_clk/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.h_flat\[134\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_427 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_65_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1058/X fanout583/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout267_A fanout267/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_1193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_942 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[22\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout434_A fanout443/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[21\]_sky130_fd_sc_hd__mux2_1_A1_S fanout220/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold930/A fanout50/X fanout79/X hold1179/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[2\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X m_blake2.m_hash256.v_q\[11\]\[0\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[25\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ sky130_fd_sc_hd__xnor2_2
XTAP_TAPCELL_ROW_46_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[247\]_sky130_fd_sc_hd__nor2_2_B/Y m_blake2.m_hash256.v_q\[7\]\[23\]_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[255\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_52_1355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_fanout222_X fanout222/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[0\]\[2\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR VPWR
+ hold655/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_59_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_59_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold350 hold350/A VGND VGND VPWR VPWR hold350/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold361 hold361/A VGND VGND VPWR VPWR hold361/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 hold372/A VGND VGND VPWR VPWR hold372/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 hold383/A VGND VGND VPWR VPWR hold383/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 hold394/A VGND VGND VPWR VPWR hold394/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_A1
+ fanout301/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[18\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout285/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout146/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A fanout83/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__and3b_2_A_N
+ m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand3_2_C/B
+ sky130_fd_sc_hd__and3b_1
XTAP_TAPCELL_ROW_5_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X_X m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.v_q\[15\]\[3\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[3\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A/X
+ sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.m_matrix\[3\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold762/X m_blake2.m_hash256.m_matrix\[4\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout555/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[3\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1050 hold1050/A VGND VGND VPWR VPWR hold1050/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[209\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xhold1072 hold1072/A VGND VGND VPWR VPWR hold1072/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2_A2 m_io.m_config.ll_q\[18\]_sky130_fd_sc_hd__o221a_2_B2/A2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1061 hold1061/A VGND VGND VPWR VPWR hold1061/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1083 hold1083/A VGND VGND VPWR VPWR hold1083/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR fanout477/A sky130_fd_sc_hd__dfxtp_1
Xhold1094 hold1094/A VGND VGND VPWR VPWR hold1094/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__a221o_2_A1 hold534/A fanout276/X
+ m_blake2.m_hash256.v_q\[14\]\[12\]_sky130_fd_sc_hd__or2_2_A/X fanout186/X fanout272/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__a221o_2_A1/X
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_43_clk/X
+ m_blake2.m_hash256.h_flat\[175\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold181/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout231/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_16_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[9\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y
+ hold1254/A m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__and3_2_B/C
+ fanout421/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[50\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X/B1
+ sky130_fd_sc_hd__a21oi_1
Xm_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[184\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold128/X fanout321/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[176\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y
+ fanout288/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_39_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__nand2_2_A_A m_blake2.m_hash256.g_b\[29\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_876 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_898 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B fanout429/X hold182/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[80\]_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_3_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D
+ m_blake2.m_hash256.m_g.a_q\[12\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[13\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[14\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D/Y
+ sky130_fd_sc_hd__nor4_2
Xm_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__or2_2_A hold360/A fanout246/X VGND VGND
+ VPWR VPWR m_io.m_config.ll_q\[45\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__mux2_1_A0 hold310/A m_blake2.m_hash256.h_flat\[197\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout397/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[5\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_64_1259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A
+ m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A/Y m_blake2.m_hash256.m_g.m_add_1.x2_i\[11\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[11\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_4
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout136/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__and2_2_B fanout440/X hold27/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[151\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
XFILLER_77_894 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_B1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_717 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2
+ fanout278/X m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[57\]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2/Y
+ fanout346/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[89\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2/X
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__a21o_2_A1/B1 m_blake2.m_hash256.m_g.m_add_1.x2_i\[21\]_sky130_fd_sc_hd__nor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/B
+ sky130_fd_sc_hd__nor2_1
XFILLER_45_780 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A0 hold228/A m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout522/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[182\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X_sky130_fd_sc_hd__xnor2_2_B_A
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[10\]\[13\]_sky130_fd_sc_hd__mux2_1_A0 hold742/X m_blake2.m_hash256.v_q\[9\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout236/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X
+ fanout257/X m_blake2.m_hash256.v_q\[6\]\[20\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X/B1
+ fanout395/X fanout179/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/A2
+ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_41_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_41_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q m_blake2.m_hash256.m_matrix\[1\]\[22\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ fanout569/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_670 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A/Y
+ m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A/B
+ m_blake2.m_hash256.m_g.b_q\[18\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.b_q\[19\]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[16\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A/X
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__xnor2_2_A hold694/A hold392/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__a22o_2_A1 hold592/A fanout188/X
+ fanout195/X hold645/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[0\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_8_clk clkload0/A VGND VGND VPWR VPWR clkbuf_leaf_8_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[1\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_54_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.m_g.d_q\[11\]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X
+ m_blake2.m_hash256.v_q\[15\]\[19\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xfanout104 fanout107/A VGND VGND VPWR VPWR fanout104/X sky130_fd_sc_hd__buf_4
Xfanout115 fanout115/A VGND VGND VPWR VPWR fanout115/X sky130_fd_sc_hd__clkbuf_2
Xfanout126 fanout127/A VGND VGND VPWR VPWR fanout126/X sky130_fd_sc_hd__clkbuf_4
Xfanout137 fanout139/X VGND VGND VPWR VPWR fanout137/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__a22o_2_A1 hold507/A fanout192/X
+ fanout200/X hold824/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[12\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout384_A fanout385/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout159 fanout160/X VGND VGND VPWR VPWR fanout159/X sky130_fd_sc_hd__buf_4
Xfanout148 fanout151/X VGND VGND VPWR VPWR fanout148/X sky130_fd_sc_hd__clkbuf_4
XFILLER_41_1023 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.m_matrix\[10\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[10\]\[13\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1025/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X
+ hold706/A fanout66/X fanout38/X hold1211/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X/C1
+ sky130_fd_sc_hd__a22o_1
XFILLER_27_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[12\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_A2
+ fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_769 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout172_X fanout172/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_2_0_clk clkbuf_0_clk/X VGND VGND VPWR VPWR clkbuf_3_2_0_clk/X sky130_fd_sc_hd__clkbuf_8
Xm_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1/Y
+ m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[11\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ sky130_fd_sc_hd__nor2_2
XFILLER_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_920 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_964 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout437_X fanout437/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[5\]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_B
+ fanout249/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/A m_blake2.m_hash256.v_q\[12\]\[21\]_sky130_fd_sc_hd__a221o_2_A1/B2
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__o21ai_2_A1/A2
+ sky130_fd_sc_hd__and3_1
Xdata\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_20_clk/X data\[0\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_1114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.v_q\[15\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/A1 fanout210/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[14\]\[15\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xdata\[1\]_sky130_fd_sc_hd__mux2_1_A1 hold14/X hold12/X fanout589/X VGND VGND VPWR
+ VPWR data\[1\]_sky130_fd_sc_hd__mux2_1_A1/X sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[14\]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1
+ fanout240/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_73_clk/X
+ m_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR m_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[28\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout198/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.d_q\[24\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkbuf_leaf_48_clk/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_9_clk/X
+ m_blake2.m_hash256.v_q\[11\]\[10\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold908/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0 hold314/A m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout378/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[1\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold180 hold180/A VGND VGND VPWR VPWR hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A1
+ m_blake2.m_hash256.m_g.a0\[7\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X/A3
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[6\]_sky130_fd_sc_hd__xor2_2_X/B sky130_fd_sc_hd__nand2_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold191 hold191/A VGND VGND VPWR VPWR hold191/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[11\]\[11\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[9\]\[11\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold695/X fanout220/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[11\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_809 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[7\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[7\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[6\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1243/X m_blake2.m_hash256.m_matrix\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout576/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[6\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_d\[18\]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B2
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_A2
+ fanout100/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_c_buf\[1\]_sky130_fd_sc_hd__o22a_2_X hold1216/A fanout175/X
+ m_blake2.m_hash256.g_c_buf\[1\]_sky130_fd_sc_hd__o22a_2_X/B1 m_blake2.m_hash256.g_c_buf\[1\]_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[1\].m_c_buf/A sky130_fd_sc_hd__o22a_1
XFILLER_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_739 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q clkload6/A m_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[13\]\[11\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[13\]\[11\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold1023/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/A
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/B
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/C
+ m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[25\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X/B2
+ sky130_fd_sc_hd__or4_1
Xm_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__mux2_1_A0 hold384/X m_blake2.m_hash256.v_q\[3\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout415/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_953 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_1063 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_B fanout288/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_912 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[36\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[9\]\[4\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[44\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/A2
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1/Y
+ sky130_fd_sc_hd__o21ai_2
Xm_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ hold1262/X fanout207/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[13\]\[12\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[28\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout116/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_967 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_70_1296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__a22o_2_A1_B1 fanout195/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/A1
+ fanout17/X m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/B1 m_blake2.m_hash256.g_y_buf\[31\]_sky130_fd_sc_hd__o22a_2_X/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[31\].m_y_buf/A sky130_fd_sc_hd__o22a_1
XFILLER_6_673 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_39_clk/X
+ m_blake2.m_hash256.v_q\[15\]\[12\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold534/A sky130_fd_sc_hd__dfxtp_1
Xm_io.m_config.ll_q\[46\]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1/B1 m_blake2.m_hash256.round_q\[0\]_sky130_fd_sc_hd__o31a_2_A1/B1
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[60\]_sky130_fd_sc_hd__a211o_2_A1/C1 sky130_fd_sc_hd__nor2_4
XFILLER_64_1089 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_1321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X
+ m_blake2.m_hash256.v_q\[1\]\[25\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold367/A sky130_fd_sc_hd__dfxtp_1
XFILLER_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_37_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_34_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[13\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold786/X hold658/X fanout580/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[13\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_886 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_867 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[230\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[7\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[238\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_43_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__and2b_2_A_N_A_N
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[16\]_sky130_fd_sc_hd__dfxtp_2_Q/Q VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_912 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[14\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold515/X m_blake2.m_hash256.m_matrix\[15\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout554/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[14\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1025/X fanout540/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[10\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B
+ m_blake2.m_hash256.m_g.a_q\[21\]_sky130_fd_sc_hd__xnor2_2_A/Y m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[20\]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B/X
+ sky130_fd_sc_hd__and2b_1
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1_A1
+ m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A
+ m_blake2.m_hash256.g_b\[30\]_sky130_fd_sc_hd__a22oi_2_B2/A1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_10_clk/X
+ m_blake2.m_hash256.v_q\[3\]\[26\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold611/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/A1
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/A2
+ m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[5\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1/X
+ sky130_fd_sc_hd__o21a_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[29\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X
+ hold813/A fanout384/X fanout194/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[4\]_sky130_fd_sc_hd__or3_2_X/B
+ sky130_fd_sc_hd__o21a_1
Xm_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A0 hold112/A m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout506/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[217\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__and2_2_B fanout433/X hold741/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__and2_2_B/X
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout599_A fanout608/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_idx_next\[1\]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_A1
+ fanout418/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.m_matrix\[2\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_CLK clkload14/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_1287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold301/A m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__and2_2_B/X fanout384/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X
+ m_blake2.m_hash256.block_idx_plus_one_q\[52\]_sky130_fd_sc_hd__and2_2_A/B fanout424/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__a31o_2_B1/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__and3b_1
Xm_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold440/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[1\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkload9/A m_blake2.m_hash256.m_matrix\[1\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold1202/A sky130_fd_sc_hd__dfxtp_1
XFILLER_70_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout45_A fanout47/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[16\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_A2
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_1345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[9\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout124/X fanout92/X
+ hold1156/A VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__mux2_1_A0 m_blake2.m_hash256.v_q\[2\]\[7\]_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.v_q\[11\]\[7\]_sky130_fd_sc_hd__mux2_1_A1/A0 fanout236/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[10\]\[7\]_sky130_fd_sc_hd__mux2_1_A0/X sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__o22a_2_A2 fanout510/X hold161/A
+ m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__o22a_2_A2/B1 m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__o22a_2_A2/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[20\]_sky130_fd_sc_hd__o22a_2_A2/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA_m_blake2.m_hash256.v_q\[10\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_S fanout235/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X
+ hold353/A fanout34/X fanout74/X hold1094/A m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[17\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X/C1
+ sky130_fd_sc_hd__a221o_1
Xm_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_60_clk/X m_blake2.m_hash256.h_flat\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold600/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload32/A m_blake2.m_hash256.v_q\[7\]\[28\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold964/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__xnor2_2_A hold796/A hold1190/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[9\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0 hold1087/X m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout153/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[9\]\[10\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_65_1343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_48_clk/X
+ m_blake2.m_hash256.m_g.a0\[27\]_sky130_fd_sc_hd__xnor2_2_Y/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_2
Xm_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ hold922/X fanout202/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[7\]\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__or2_2_B fanout498/X hold125/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[215\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_39_809 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[37\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold382/X fanout325/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[29\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/Q hold1176/X
+ fanout562/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[12\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xfanout490 fanout494/X VGND VGND VPWR VPWR fanout490/X sky130_fd_sc_hd__buf_2
Xm_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1
+ m_blake2.m_hash256.m_g.b_q\[29\]_sky130_fd_sc_hd__xor2_2_A/B m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y/B
+ m_blake2.m_hash256.m_g.b_q\[28\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[30\]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X/B1
+ sky130_fd_sc_hd__o21ai_1
XFILLER_24_1084 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1073 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_69_clk/X m_blake2.m_hash256.h_flat\[8\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold96/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_matrix\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1165/X hold880/A fanout551/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_59_1147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ hold1264/A fanout143/X fanout118/X m_blake2.m_hash256.m_matrix\[13\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[3\]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B
+ m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__nand2_2_A/Y m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[24\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nor2_2_Y
+ fanout388/X fanout253/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ sky130_fd_sc_hd__nor2_8
XFILLER_72_1314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_57_clk/X
+ m_blake2.m_hash256.v_q\[9\]\[29\]_sky130_fd_sc_hd__mux2_1_A0/X VGND VGND VPWR VPWR
+ hold674/A sky130_fd_sc_hd__dfxtp_1
XFILLER_42_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[5\]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout124/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_783 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__dfxtp_2_Q clkload23/A m_blake2.m_hash256.g_buffer\[28\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[28\]_sky130_fd_sc_hd__or2_2_A/A
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X
+ fanout255/X m_blake2.m_hash256.v_q\[6\]\[17\]_sky130_fd_sc_hd__mux2_1_A0/X m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X/B1
+ fanout367/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X/A1
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_matrix\[6\]\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold781/X hold1238/A fanout590/X VGND VGND VPWR VPWR hold782/A sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[9\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1
+ fanout46/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_764 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_742 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[15\]\[1\]_sky130_fd_sc_hd__mux2_1_A0_S fanout296/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B fanout483/X hold138/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[49\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_1077 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold927 hold927/A VGND VGND VPWR VPWR hold927/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 hold916/A VGND VGND VPWR VPWR hold916/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold905 hold905/A VGND VGND VPWR VPWR hold905/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 hold938/A VGND VGND VPWR VPWR hold938/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold949 hold949/A VGND VGND VPWR VPWR hold949/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2
+ fanout350/X m_blake2.m_hash256.v_q\[5\]\[27\]_sky130_fd_sc_hd__a22o_2_A1/X m_blake2.m_hash256.v_q\[6\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[27\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y/B1
+ sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A0 hold37/A m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout529/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_1427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_36_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[4\]\[30\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold232/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_32_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_1067 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X m_blake2.m_hash256.g_d\[9\]_sky130_fd_sc_hd__a21oi_2_Y/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.d_q\[9\]_sky130_fd_sc_hd__xor2_2_B/B
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B fanout484/X hold178/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[42\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
XFILLER_77_1203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_853 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xm_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X
+ m_blake2.m_hash256.m_matrix\[14\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q fanout89/X
+ fanout113/X m_blake2.m_hash256.m_matrix\[5\]\[15\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[15\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_38_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[9\]_sky130_fd_sc_hd__a31o_2_A3_A2 fanout476/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1/X
+ m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A/B
+ sky130_fd_sc_hd__or2_1
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout347_A fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X
+ m_io.m_config.cfg_cnt_q\[3\]_sky130_fd_sc_hd__nand3_2_C/B m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X/B
+ VGND VGND VPWR VPWR m_io.m_config.cfg_cnt_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X/C
+ sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[2\]_sky130_fd_sc_hd__mux2_1_A1_S fanout225/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2
+ fanout134/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1
+ fanout179/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_c_buf\[26\]_sky130_fd_sc_hd__a211o_2_X_A2 fanout174/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_775 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_797 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q clkload14/A m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[8\]\[10\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X
+ m_blake2.m_hash256.v_q\[6\]\[31\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold956/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_A3
+ m_blake2.m_hash256.v_q\[15\]\[13\]_sky130_fd_sc_hd__mux2_1_A0/A1 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2
+ m_blake2.m_hash256.m_g.a0\[28\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X/B2
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[26\]_sky130_fd_sc_hd__nand2_2_A/Y sky130_fd_sc_hd__nand2_1
XANTENNA_m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__mux2_1_A0_A0 m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[25\]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout66/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[12\]_sky130_fd_sc_hd__xor2_2_A/X sky130_fd_sc_hd__xor2_4
XANTENNA_fanout302_X fanout302/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1
+ fanout199/X m_blake2.m_hash256.h_flat\[237\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout192/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[173\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[20\]_sky130_fd_sc_hd__dfxtp_2_Q_D m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__o22a_2_X/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_S fanout229/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.v_q\[0\]\[21\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2
+ fanout406/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B/A
+ m_blake2.m_hash256.m_g.a_q\[4\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A/Y
+ m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B/A
+ sky130_fd_sc_hd__a21o_1
XANTENNA_m_blake2.m_hash256.g_d\[24\]_sky130_fd_sc_hd__a21oi_2_Y_A1 fanout271/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_679 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X/A1
+ m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X/A2 m_blake2.m_hash256.g_y_buf\[3\]_sky130_fd_sc_hd__o32a_2_X/A3
+ fanout19/X hold235/A VGND VGND VPWR VPWR m_blake2.m_hash256.g_buffer\[3\].m_y_buf/A
+ sky130_fd_sc_hd__o32a_1
XFILLER_21_1202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__a22o_2_A1 hold139/X fanout336/X
+ m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__a22o_2_A1/B1 fanout531/X VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[254\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__and2b_2_B m_blake2.m_hash256.m_g.b_q\[22\]_sky130_fd_sc_hd__xor2_2_A/X
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[10\]_sky130_fd_sc_hd__xnor2_2_A/A VGND VGND
+ VPWR VPWR m_blake2.m_hash256.m_g.a_q\[10\]_sky130_fd_sc_hd__a21oi_2_A1/B1 sky130_fd_sc_hd__and2b_1
XFILLER_5_1454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__a22o_2_A1 m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__nor2_2_B/B
+ fanout340/X m_blake2.m_hash256.h_flat\[141\]_sky130_fd_sc_hd__a31o_2_A3/X m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__a22o_2_A1/B2
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[133\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X
+ fanout451/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_B/X VGND VGND
+ VPWR VPWR m_blake2.m_hash256.round_q\[7\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X/A3
+ sky130_fd_sc_hd__or2_1
XFILLER_29_897 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_d\[2\]_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__o211a_2_X_B1
+ fanout237/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_856 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q clkload27/A m_blake2.m_hash256.g_b\[31\]_sky130_fd_sc_hd__xor2_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/Q
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout48_X fanout48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.m_matrix\[0\]\[1\]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_A2
+ fanout142/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[4\]_sky130_fd_sc_hd__nand2_2_A_B fanout288/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_753 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__inv_2_A
+ m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[18\]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[16\]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_A
+ fanout349/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_757 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[51\]_sky130_fd_sc_hd__dfxtp_2_Q_Q
+ m_io.m_config.ll_q\[57\]_sky130_fd_sc_hd__a221o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_974 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_72_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y_A m_blake2.m_hash256.g_b\[15\]_sky130_fd_sc_hd__inv_2_Y/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[1\]_sky130_fd_sc_hd__and4_2_B_B
+ m_io.m_config.ll_q\[7\]_sky130_fd_sc_hd__a22o_2_B2/A1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_948 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.m_g.a0\[0\]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_X
+ m_blake2.m_hash256.m_matrix\[0\]\[0\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__xnor2_2_A hold313/A hold672/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[0\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_1
XFILLER_74_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_1133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X m_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[6\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_io.m_config.kk_q\[4\]_sky130_fd_sc_hd__or2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_1231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_1177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_34_clk/X
+ m_blake2.m_hash256.h_flat\[243\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold741/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_61_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__dfxtp_2_Q clkload17/A m_blake2.m_hash256.h_flat\[122\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold212/A sky130_fd_sc_hd__dfxtp_1
Xhold702 hold702/A VGND VGND VPWR VPWR hold702/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 hold713/A VGND VGND VPWR VPWR hold713/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold746 hold746/A VGND VGND VPWR VPWR hold746/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 hold724/A VGND VGND VPWR VPWR hold724/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold735 hold735/A VGND VGND VPWR VPWR hold735/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[252\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold265/X fanout336/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[244\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xhold757 hold757/A VGND VGND VPWR VPWR hold757/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold779 hold779/A VGND VGND VPWR VPWR hold779/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 hold768/A VGND VGND VPWR VPWR hold768/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_S fanout157/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[185\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[5\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[193\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XFILLER_44_1213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xm_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[131\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold56/X fanout334/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[123\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout297_A fanout299/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[22\]_sky130_fd_sc_hd__mux2_1_A0_S fanout302/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_1257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__a22o_2_A1 hold344/A fanout290/X
+ fanout284/X hold754/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[1\]\[2\]_sky130_fd_sc_hd__a22o_2_A1/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_73_907 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X
+ hold251/A m_blake2.m_hash256.h_flat\[147\]_sky130_fd_sc_hd__or2_2_B/X fanout375/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X/B1 sky130_fd_sc_hd__mux2_1
XFILLER_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1011 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_fanout464_A fanout465/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[15\]_sky130_fd_sc_hd__o22a_2_A1_B1 fanout172/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o311a_2_X
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X/A
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X/A ANTENNA_6/DIODE m_blake2.m_hash256.g_b\[12\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2/X
+ m_blake2.m_hash256.m_g.a0\[12\]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a0\[14\]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_80_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout252_X fanout252/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_1028 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_m_blake2.m_hash256.g_c_buf\[3\]_sky130_fd_sc_hd__a21o_2_X_A1 m_blake2.m_hash256.g_c_buf\[7\]_sky130_fd_sc_hd__a21o_2_X/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1
+ fanout290/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.h_flat\[32\]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_B2
+ fanout278/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_68_clk/X m_blake2.m_hash256.g_buffer\[0\].m_c_buf/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.c_q\[0\]_sky130_fd_sc_hd__or2_2_A/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1/B2 m_blake2.m_hash256.block_idx_plus_one_q\[4\]_sky130_fd_sc_hd__and4_2_C/D
+ fanout427/X VGND VGND VPWR VPWR m_blake2.m_hash256.block_idx_plus_one_q\[2\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
Xm_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B/A
+ hold1014/A VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[18\]_sky130_fd_sc_hd__xnor2_2_B/Y
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_matrix\[2\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1229/X hold1003/X fanout557/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[28\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.v_q\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ m_blake2.m_hash256.v_q\[11\]\[5\]_sky130_fd_sc_hd__mux2_1_A1/A0 hold844/X fanout223/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[8\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__dfxtp_2_Q_Q m_blake2.m_hash256.m_g.m_add_1.x2_i\[4\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_716 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__mux2_1_A0 hold437/A m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout513/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[250\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_749 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_49_1157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold366/X m_blake2.m_hash256.v_q\[7\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X/A0
+ fanout157/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[1\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A/A
+ fanout487/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[128\]_sky130_fd_sc_hd__nor2_2_A/Y
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S
+ fanout159/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/A
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.a_q\[24\]_sky130_fd_sc_hd__or2_2_A/X sky130_fd_sc_hd__or2_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[11\]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y
+ m_blake2.m_hash256.g_b\[11\]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.block_idx_plus_one_q\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_A2
+ m_blake2.m_hash256.block_idx_plus_one_q\[16\]_sky130_fd_sc_hd__and4_2_C/D VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_1 hold293/A m_blake2.m_hash256.h_flat\[138\]_sky130_fd_sc_hd__and2_2_B/X
+ fanout370/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[10\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__xnor2_2_A hold458/A hold1230/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[23\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold62 hold62/A VGND VGND VPWR VPWR hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A VGND VGND VPWR VPWR hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A VGND VGND VPWR VPWR hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A VGND VGND VPWR VPWR hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_A
+ m_blake2.m_hash256.m_g.m_add_1.x2_i\[25\]_sky130_fd_sc_hd__inv_2_A/Y VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_matrix\[9\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold353/X hold369/X fanout580/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[9\]\[17\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_3_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[11\]\[1\]_sky130_fd_sc_hd__o22a_2_A1_B1 fanout171/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_38_clk/X
+ m_blake2.m_hash256.h_flat\[148\]_sky130_fd_sc_hd__mux2_1_A1/X VGND VGND VPWR VPWR
+ hold26/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_A1 hash\[0\]_sky130_fd_sc_hd__or2_2_B/B
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1211/X hold1183/X fanout580/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[9\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_14_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/B m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/C
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.b_q\[14\]_sky130_fd_sc_hd__nand3_2_A/Y
+ sky130_fd_sc_hd__nand3_2
XFILLER_34_1459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[157\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold90/X fanout339/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[149\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_61_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_74_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[8\]_sky130_fd_sc_hd__a32o_2_A1_A3 fanout250/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_58_clk/X m_blake2.m_hash256.h_flat\[61\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold152/A sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_74_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_4 ANTENNA_4/DIODE VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.m_matrix\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold1101/X hold920/X fanout542/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[2\]\[5\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X
+ fanout237/X m_blake2.m_hash256.v_q\[13\]\[0\]_sky130_fd_sc_hd__a221o_2_A1/X fanout270/X
+ m_io.m_config.ll_q\[0\]_sky130_fd_sc_hd__o2bb2a_2_A1_N/X VGND VGND VPWR VPWR m_blake2.m_hash256.g_d\[0\]_sky130_fd_sc_hd__or3_2_X/C
+ sky130_fd_sc_hd__a22o_1
Xm_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[70\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold50/X fanout331/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[62\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[7\]\[17\]_sky130_fd_sc_hd__mux2_1_A1/A0
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[2\]\[23\]_sky130_fd_sc_hd__mux2_1_A0_S fanout415/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_1457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_67_734 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1037 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_745 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_6_clk_A clkbuf_3_0_0_clk/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_io.m_config.ll_q\[37\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2
+ fanout168/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__xnor2_2_A hold283/A hold1163/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[25\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_50_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_981 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_1_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.m_matrix\[0\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold852/X hold675/X fanout571/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[0\]\[14\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_78_1342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__and2_2_B fanout432/X hold36/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[154\]_sky130_fd_sc_hd__and2_2_B/X sky130_fd_sc_hd__and2_1
Xm_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y
+ fanout474/X m_blake2.m_hash256.g_idx_next\[2\]_sky130_fd_sc_hd__o21ai_2_A1/Y fanout481/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_idx_q\[0\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y/B
+ sky130_fd_sc_hd__o21ai_1
XFILLER_23_815 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_63_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_m_blake2.m_hash256.v_q\[12\]\[8\]_sky130_fd_sc_hd__a221o_2_A1_C1 fanout268/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_m_blake2.m_hash256.v_q\[1\]\[13\]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1
+ fanout104/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_63_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2_A2 fanout265/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_42_clk/X m_io.m_config.ll_q\[54\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold240/A sky130_fd_sc_hd__dfxtp_1
XFILLER_50_678 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A0 hold100/A m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout515/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[155\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_30_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q clkload25/A m_blake2.m_hash256.v_q\[8\]\[3\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hold775/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_D_sky130_fd_sc_hd__o311a_2_X
+ fanout455/X m_blake2.m_hash256.round_q\[9\]_sky130_fd_sc_hd__or2_2_A/X m_blake2.m_hash256.round_q\[8\]_sky130_fd_sc_hd__or2_2_A/X
+ fanout401/X fanout468/X VGND VGND VPWR VPWR m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C/D
+ sky130_fd_sc_hd__o311a_1
Xhold510 hold510/A VGND VGND VPWR VPWR hold510/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__xnor2_2_A hold347/A hold519/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[6\]\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
Xhold532 hold532/A VGND VGND VPWR VPWR hold532/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 hold521/A VGND VGND VPWR VPWR hold521/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 hold554/A VGND VGND VPWR VPWR hold554/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 hold543/A VGND VGND VPWR VPWR hold543/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_11_1289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_57_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold587 hold587/A VGND VGND VPWR VPWR hold587/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 hold576/A VGND VGND VPWR VPWR hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 hold565/A VGND VGND VPWR VPWR hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 hold598/A VGND VGND VPWR VPWR hold598/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1 hold242/A m_blake2.m_hash256.h_flat\[171\]_sky130_fd_sc_hd__or2_2_B/X
+ fanout377/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[5\]\[11\]_sky130_fd_sc_hd__mux2_1_A0_1/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_y_buf\[11\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1221 hold1221/A VGND VGND VPWR VPWR hold1221/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1210 hold1210/A VGND VGND VPWR VPWR hold1210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1232 hold1232/A VGND VGND VPWR VPWR hold1232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1243 hold1243/A VGND VGND VPWR VPWR hold1243/X sky130_fd_sc_hd__dlygate4sd3_1
Xm_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B fanout496/X hold88/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[39\]_sky130_fd_sc_hd__or2_2_B/X sky130_fd_sc_hd__or2_1
Xm_blake2.m_hash256.v_q\[14\]\[4\]_sky130_fd_sc_hd__dfxtp_2_Q clkload33/A m_blake2.m_hash256.v_q\[14\]\[4\]_sky130_fd_sc_hd__mux2_1_A0/X
+ VGND VGND VPWR VPWR hold457/A sky130_fd_sc_hd__dfxtp_1
Xhold1254 hold1254/A VGND VGND VPWR VPWR hold1254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold1265 hold1265/A VGND VGND VPWR VPWR hold1265/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_m_blake2.m_hash256.h_flat\[33\]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1
+ fanout289/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_1426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_m_blake2.m_hash256.g_y_buf\[4\]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1
+ fanout72/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X
+ hold361/A fanout80/X fanout64/X hold1113/A m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X/C1
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_y_buf\[21\]_sky130_fd_sc_hd__o32a_2_X/A3
+ sky130_fd_sc_hd__a221o_1
XPHY_EDGE_ROW_11_Left_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__xnor2_2_A hold444/A hold1194/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[4\]\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XFILLER_40_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xm_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1
+ m_blake2.m_hash256.m_g.c_q\[12\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.c_q\[11\]_sky130_fd_sc_hd__a21oi_2_A1/Y m_blake2.m_hash256.m_g.c_q\[13\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B/X
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1/Y VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.c_q\[15\]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1/X
+ sky130_fd_sc_hd__o41a_1
XTAP_TAPCELL_ROW_24_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_56_clk/X m_blake2.m_hash256.h_flat\[87\]_sky130_fd_sc_hd__mux2_1_A1/X
+ VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/A
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/B VGND VGND VPWR VPWR
+ m_blake2.m_hash256.m_g.b_q\[26\]_sky130_fd_sc_hd__xnor2_2_A/Y sky130_fd_sc_hd__xnor2_4
Xm_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[27\]_sky130_fd_sc_hd__or2_2_B/X m_blake2.m_hash256.v_q\[0\]\[27\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[35\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
Xm_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A
+ m_blake2.m_hash256.m_g.b_q\[5\]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B/Y
+ m_blake2.m_hash256.m_g.a_q\[27\]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[24\]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2/B1
+ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_24_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_m_blake2.m_hash256.v_q\[14\]\[19\]_sky130_fd_sc_hd__mux2_1_A0_S fanout209/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__xnor2_2_A m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__o22a_2_X/X
+ m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__and2_2_A/B VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[1\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__a221oi_2_A1_A1 m_blake2.m_hash256.m_g.c_q\[3\]_sky130_fd_sc_hd__xnor2_2_A/A
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__mux2_1_A0 hold619/A m_io.m_config.kk_q\[0\]_sky130_fd_sc_hd__mux2_1_A1/X
+ fanout366/X VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[0\]\[8\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_9_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.g_b\[6\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1
+ fanout180/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A1 m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__mux2_1_A0/X
+ hold1102/X fanout318/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[88\]_sky130_fd_sc_hd__mux2_1_A1/X
+ sky130_fd_sc_hd__mux2_1
Xm_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/A
+ m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y/B
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[20\]_sky130_fd_sc_hd__nor2_2_A/B sky130_fd_sc_hd__xnor2_1
XFILLER_16_1189 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_blake2.m_hash256.m_matrix\[5\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X
+ hold736/X hold414/X fanout572/X VGND VGND VPWR VPWR m_blake2.m_hash256.m_matrix\[5\]\[23\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhash\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkload28/A hash\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D
+ VGND VGND VPWR VPWR hash\[6\]_sky130_fd_sc_hd__or2_2_B/B sky130_fd_sc_hd__dfxtp_4
XANTENNA_m_blake2.m_hash256.v_q\[6\]\[13\]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_A1
+ fanout257/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xm_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X
+ hold259/X fanout165/X m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__or2_2_A/X fanout619/X
+ VGND VGND VPWR VPWR m_io.m_config.ll_q\[31\]_sky130_fd_sc_hd__dfxtp_2_Q/D sky130_fd_sc_hd__o211a_1
XANTENNA_m_blake2.m_hash256.v_q\[3\]\[24\]_sky130_fd_sc_hd__mux2_1_A0_S fanout418/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_1143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nand4_2_C
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1/X
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2/B
+ m_blake2.m_hash256.round_q\[5\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B/Y
+ m_blake2.m_hash256.round_q\[1\]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B/Y
+ VGND VGND VPWR VPWR fanout103/A sky130_fd_sc_hd__nand4_1
Xm_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B fanout494/X hold261/A VGND
+ VGND VPWR VPWR m_blake2.m_hash256.h_flat\[93\]_sky130_fd_sc_hd__nor2_2_B/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_1285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_m_blake2.m_hash256.g_b\[19\]_sky130_fd_sc_hd__o22a_2_X_B2 fanout181/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xm_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X
+ fanout345/X m_blake2.m_hash256.v_q\[5\]\[17\]_sky130_fd_sc_hd__a22o_2_A1/X fanout177/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.g_b\[17\]_sky130_fd_sc_hd__o22a_2_X/A2 sky130_fd_sc_hd__a21o_1
Xm_blake2.m_hash256.m_matrix\[14\]\[8\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_15_clk/X
+ hold1059/X VGND VGND VPWR VPWR hold1058/A sky130_fd_sc_hd__dfxtp_1
XFILLER_45_951 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/A
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.m_add_1.x2_i\[14\]_sky130_fd_sc_hd__inv_2_A/Y
+ sky130_fd_sc_hd__clkinv_2
XFILLER_16_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xm_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__a211o_2_A1 m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__xor2_2_B/B
+ fanout282/X m_blake2.m_hash256.v_q\[1\]\[14\]_sky130_fd_sc_hd__a22o_2_A1/X fanout386/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.v_q\[2\]\[14\]_sky130_fd_sc_hd__a211o_2_A1/X
+ sky130_fd_sc_hd__a211o_1
Xm_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A0 hold71/A m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ fanout525/X VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[94\]_sky130_fd_sc_hd__mux2_1_A0/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_13_870 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.h_flat\[96\]_sky130_fd_sc_hd__and2_2_B_A fanout429/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xm_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_47_clk/X
+ m_blake2.m_hash256.block_idx_plus_one_q\[42\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND
+ VGND VPWR VPWR m_io.m_config.ll_q\[48\]_sky130_fd_sc_hd__a22oi_2_B2/A1 sky130_fd_sc_hd__dfxtp_1
Xm_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_28_clk/X m_blake2.m_hash256.m_g.a0\[1\]_sky130_fd_sc_hd__and2b_2_X/X
+ VGND VGND VPWR VPWR m_blake2.m_hash256.m_g.a_q\[1\]_sky130_fd_sc_hd__inv_2_A/A sky130_fd_sc_hd__dfxtp_1
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xm_blake2.m_hash256.m_matrix\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q clkbuf_leaf_72_clk/X
+ m_blake2.m_hash256.m_matrix\[9\]\[6\]_sky130_fd_sc_hd__dfxtp_2_Q/D VGND VGND VPWR
+ VPWR hold1049/A sky130_fd_sc_hd__dfxtp_1
XFILLER_67_1032 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0_A1 m_blake2.m_hash256.v_q\[9\]\[27\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout319 fanout320/X VGND VGND VPWR VPWR fanout319/X sky130_fd_sc_hd__clkbuf_4
Xfanout308 fanout308/A VGND VGND VPWR VPWR fanout308/X sky130_fd_sc_hd__clkbuf_4
XFILLER_59_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xm_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B
+ m_blake2.m_hash256.h_flat\[198\]_sky130_fd_sc_hd__and2_2_B/X m_blake2.m_hash256.v_q\[6\]\[6\]_sky130_fd_sc_hd__xnor2_2_A/Y
+ VGND VGND VPWR VPWR m_blake2.m_hash256.h_flat\[206\]_sky130_fd_sc_hd__mux2_1_A0/A1
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X_B1 m_blake2.m_hash256.g_c_buf\[31\]_sky130_fd_sc_hd__a221o_2_X/B1
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
.ends

