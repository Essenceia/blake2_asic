module tt_um_essen (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire block_first;
 wire block_first_sky130_fd_sc_hd__a32o_2_B2_A1;
 wire block_first_sky130_fd_sc_hd__dfxtp_2_Q_D;
 wire block_first_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B;
 wire block_last;
 wire block_last_sky130_fd_sc_hd__a22o_2_B2_A2;
 wire block_last_sky130_fd_sc_hd__a22o_2_B2_B1;
 wire block_last_sky130_fd_sc_hd__dfxtp_2_Q_D;
 wire block_last_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B;
 wire \data[0] ;
 wire \data[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data[1] ;
 wire \data[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data[2] ;
 wire \data[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data[3] ;
 wire \data[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data[4] ;
 wire \data[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data[5] ;
 wire \data[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data[6] ;
 wire \data[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data[7] ;
 wire \data[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \data_idx[0] ;
 wire \data_idx[0]_sky130_fd_sc_hd__and4_2_B_X ;
 wire \data_idx[1] ;
 wire \data_idx[2] ;
 wire \data_idx[3] ;
 wire \data_idx[3]_sky130_fd_sc_hd__and4_2_A_X ;
 wire \data_idx[4] ;
 wire \data_idx[5] ;
 wire data_v;
 wire ena_sky130_fd_sc_hd__or2_2_B_A;
 wire \hash[0] ;
 wire \hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \hash[0]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \hash[0]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ;
 wire \hash[1] ;
 wire \hash[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \hash[1]_sky130_fd_sc_hd__mux2_1_A1_X ;
 wire \hash[2] ;
 wire \hash[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \hash[2]_sky130_fd_sc_hd__mux2_1_A1_X ;
 wire \hash[2]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2_Y ;
 wire \hash[3] ;
 wire \hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \hash[4] ;
 wire \hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \hash[4]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \hash[5] ;
 wire \hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ;
 wire \hash[6] ;
 wire \hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \hash[6]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \hash[7] ;
 wire \hash[7]_sky130_fd_sc_hd__and2_2_B_A ;
 wire \hash[7]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire hash_v;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[0] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[10] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[11] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[12] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[13] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[14] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[15] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[16] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[17] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[18] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[19] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[1] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[20] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[21] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[22] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[23] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[24] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[25] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[26] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[27] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[28] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[29] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[2] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[30] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[31] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[32] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[33] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[34] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[35] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[36] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[37] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[38] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[39] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[3] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[40] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[41] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[42] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[43] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[44] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[45] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[46] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[47] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[48] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[49] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[4] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[50] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[51] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[52] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[53] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[54] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[55] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[56] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[57] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[5] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[6] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[7] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_A2 ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[8] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[9] ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.f_finished ;
 wire \m_blake2.m_hash256.f_finished_q ;
 wire \m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_A ;
 wire \m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.first_block_q ;
 wire \m_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.fsm_q[0] ;
 wire \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.fsm_q[1] ;
 wire \m_blake2.m_hash256.fsm_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.fsm_q[2] ;
 wire \m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X_B1 ;
 wire \m_blake2.m_hash256.fsm_q[3] ;
 wire \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2 ;
 wire \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1 ;
 wire \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.fsm_q[4] ;
 wire \m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2 ;
 wire \m_blake2.m_hash256.fsm_q[5] ;
 wire \m_blake2.m_hash256.fsm_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.g_b[0] ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[10] ;
 wire \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[11] ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[12] ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.g_b[13] ;
 wire \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[14] ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.g_b[15] ;
 wire \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[16] ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[17] ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.g_b[18] ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_A ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.g_b[19] ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_X ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a221o_2_C1_X ;
 wire \m_blake2.m_hash256.g_b[1] ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[20] ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_Y ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2_Y ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[21] ;
 wire \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[22] ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.g_b[23] ;
 wire \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[24] ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[25] ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[26] ;
 wire \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[27] ;
 wire \m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[28] ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[29] ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.g_b[2] ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A1_N ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A2_N ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_X ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[30] ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A2 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_Y ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[31] ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[3] ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_A2 ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_X ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[4] ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[5] ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[6] ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_b[7] ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[8] ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_Y ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.g_b[9] ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ;
 wire \m_blake2.m_hash256.g_c[0] ;
 wire \m_blake2.m_hash256.g_c[10] ;
 wire \m_blake2.m_hash256.g_c[11] ;
 wire \m_blake2.m_hash256.g_c[12] ;
 wire \m_blake2.m_hash256.g_c[13] ;
 wire \m_blake2.m_hash256.g_c[14] ;
 wire \m_blake2.m_hash256.g_c[15] ;
 wire \m_blake2.m_hash256.g_c[16] ;
 wire \m_blake2.m_hash256.g_c[17] ;
 wire \m_blake2.m_hash256.g_c[18] ;
 wire \m_blake2.m_hash256.g_c[19] ;
 wire \m_blake2.m_hash256.g_c[1] ;
 wire \m_blake2.m_hash256.g_c[20] ;
 wire \m_blake2.m_hash256.g_c[21] ;
 wire \m_blake2.m_hash256.g_c[22] ;
 wire \m_blake2.m_hash256.g_c[23] ;
 wire \m_blake2.m_hash256.g_c[24] ;
 wire \m_blake2.m_hash256.g_c[25] ;
 wire \m_blake2.m_hash256.g_c[26] ;
 wire \m_blake2.m_hash256.g_c[27] ;
 wire \m_blake2.m_hash256.g_c[28] ;
 wire \m_blake2.m_hash256.g_c[29] ;
 wire \m_blake2.m_hash256.g_c[2] ;
 wire \m_blake2.m_hash256.g_c[30] ;
 wire \m_blake2.m_hash256.g_c[31] ;
 wire \m_blake2.m_hash256.g_c[3] ;
 wire \m_blake2.m_hash256.g_c[4] ;
 wire \m_blake2.m_hash256.g_c[5] ;
 wire \m_blake2.m_hash256.g_c[6] ;
 wire \m_blake2.m_hash256.g_c[7] ;
 wire \m_blake2.m_hash256.g_c[8] ;
 wire \m_blake2.m_hash256.g_c[9] ;
 wire \m_blake2.m_hash256.g_c_buf[0] ;
 wire \m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[10] ;
 wire \m_blake2.m_hash256.g_c_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[11] ;
 wire \m_blake2.m_hash256.g_c_buf[11]_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[12] ;
 wire \m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[13] ;
 wire \m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_c_buf[14] ;
 wire \m_blake2.m_hash256.g_c_buf[14]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[15] ;
 wire \m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_c_buf[16] ;
 wire \m_blake2.m_hash256.g_c_buf[16]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[17] ;
 wire \m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_D1 ;
 wire \m_blake2.m_hash256.g_c_buf[18] ;
 wire \m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_D1 ;
 wire \m_blake2.m_hash256.g_c_buf[19] ;
 wire \m_blake2.m_hash256.g_c_buf[19]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[1] ;
 wire \m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_c_buf[20] ;
 wire \m_blake2.m_hash256.g_c_buf[20]_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_c_buf[21] ;
 wire \m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[22] ;
 wire \m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_D1 ;
 wire \m_blake2.m_hash256.g_c_buf[23] ;
 wire \m_blake2.m_hash256.g_c_buf[23]_sky130_fd_sc_hd__o311a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[24] ;
 wire \m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[25] ;
 wire \m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_B2 ;
 wire \m_blake2.m_hash256.g_c_buf[26] ;
 wire \m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[27] ;
 wire \m_blake2.m_hash256.g_c_buf[27]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[27]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_c_buf[28] ;
 wire \m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[29] ;
 wire \m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_c_buf[2] ;
 wire \m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[30] ;
 wire \m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[31] ;
 wire \m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[3] ;
 wire \m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ;
 wire \m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[4] ;
 wire \m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[5] ;
 wire \m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_c_buf[6] ;
 wire \m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[7] ;
 wire \m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[8] ;
 wire \m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_c_buf[9] ;
 wire \m_blake2.m_hash256.g_c_buf[9]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[0] ;
 wire \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_A ;
 wire \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_B ;
 wire \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C ;
 wire \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B2 ;
 wire \m_blake2.m_hash256.g_d[10] ;
 wire \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[11] ;
 wire \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A1 ;
 wire \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[12] ;
 wire \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[13] ;
 wire \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2 ;
 wire \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[14] ;
 wire \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ;
 wire \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ;
 wire \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ;
 wire \m_blake2.m_hash256.g_d[15] ;
 wire \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[16] ;
 wire \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[17] ;
 wire \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[18] ;
 wire \m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_A2_N ;
 wire \m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_d[19] ;
 wire \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[1] ;
 wire \m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[20] ;
 wire \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[21] ;
 wire \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[22] ;
 wire \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[23] ;
 wire \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[24] ;
 wire \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ;
 wire \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ;
 wire \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ;
 wire \m_blake2.m_hash256.g_d[25] ;
 wire \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A1 ;
 wire \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[26] ;
 wire \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[27] ;
 wire \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A1 ;
 wire \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[28] ;
 wire \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ;
 wire \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ;
 wire \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ;
 wire \m_blake2.m_hash256.g_d[29] ;
 wire \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[2] ;
 wire \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__o211a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1 ;
 wire \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__o221a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_d[30] ;
 wire \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[31] ;
 wire \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2 ;
 wire \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[3] ;
 wire \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__o211a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_d[4] ;
 wire \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_A ;
 wire \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_B ;
 wire \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C ;
 wire \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[5] ;
 wire \m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[6] ;
 wire \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[7] ;
 wire \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[8] ;
 wire \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[9] ;
 wire \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ;
 wire \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_idx_next[0] ;
 wire \m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.g_idx_next[1] ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ;
 wire \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X ;
 wire \m_blake2.m_hash256.g_idx_next[2] ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_1_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_1_Y ;
 wire \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.g_idx_q[0] ;
 wire \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.g_idx_q[1] ;
 wire \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.g_idx_q[2] ;
 wire \m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C ;
 wire \m_blake2.m_hash256.g_y[0] ;
 wire \m_blake2.m_hash256.g_y[10] ;
 wire \m_blake2.m_hash256.g_y[11] ;
 wire \m_blake2.m_hash256.g_y[12] ;
 wire \m_blake2.m_hash256.g_y[13] ;
 wire \m_blake2.m_hash256.g_y[14] ;
 wire \m_blake2.m_hash256.g_y[15] ;
 wire \m_blake2.m_hash256.g_y[16] ;
 wire \m_blake2.m_hash256.g_y[17] ;
 wire \m_blake2.m_hash256.g_y[18] ;
 wire \m_blake2.m_hash256.g_y[19] ;
 wire \m_blake2.m_hash256.g_y[1] ;
 wire \m_blake2.m_hash256.g_y[20] ;
 wire \m_blake2.m_hash256.g_y[21] ;
 wire \m_blake2.m_hash256.g_y[22] ;
 wire \m_blake2.m_hash256.g_y[23] ;
 wire \m_blake2.m_hash256.g_y[24] ;
 wire \m_blake2.m_hash256.g_y[25] ;
 wire \m_blake2.m_hash256.g_y[26] ;
 wire \m_blake2.m_hash256.g_y[27] ;
 wire \m_blake2.m_hash256.g_y[28] ;
 wire \m_blake2.m_hash256.g_y[29] ;
 wire \m_blake2.m_hash256.g_y[2] ;
 wire \m_blake2.m_hash256.g_y[30] ;
 wire \m_blake2.m_hash256.g_y[31] ;
 wire \m_blake2.m_hash256.g_y[3] ;
 wire \m_blake2.m_hash256.g_y[4] ;
 wire \m_blake2.m_hash256.g_y[5] ;
 wire \m_blake2.m_hash256.g_y[6] ;
 wire \m_blake2.m_hash256.g_y[7] ;
 wire \m_blake2.m_hash256.g_y[8] ;
 wire \m_blake2.m_hash256.g_y[9] ;
 wire \m_blake2.m_hash256.g_y_buf[0] ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[10] ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_y_buf[11] ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[12] ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[13] ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[14] ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[15] ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_y_buf[16] ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[17] ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[18] ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[19] ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[1] ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[20] ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[21] ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[22] ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[23] ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[24] ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[25] ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_y_buf[26] ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_y_buf[27] ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[28] ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[29] ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[2] ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_y_buf[30] ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[31] ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[3] ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[4] ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[5] ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.g_y_buf[6] ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[7] ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[8] ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[9] ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.h_flat[100] ;
 wire \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[101] ;
 wire \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[102] ;
 wire \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[103] ;
 wire \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[104] ;
 wire \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[105] ;
 wire \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[106] ;
 wire \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[107] ;
 wire \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[108] ;
 wire \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[109] ;
 wire \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[10] ;
 wire \m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[110] ;
 wire \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[111] ;
 wire \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[112] ;
 wire \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[113] ;
 wire \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[114] ;
 wire \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[115] ;
 wire \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[116] ;
 wire \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[117] ;
 wire \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[118] ;
 wire \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[119] ;
 wire \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[11] ;
 wire \m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2_B1 ;
 wire \m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2_B2 ;
 wire \m_blake2.m_hash256.h_flat[120] ;
 wire \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[121] ;
 wire \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[122] ;
 wire \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[123] ;
 wire \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[124] ;
 wire \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[125] ;
 wire \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[126] ;
 wire \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[127] ;
 wire \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[128] ;
 wire \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[129] ;
 wire \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[12] ;
 wire \m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2_B1 ;
 wire \m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2_B2 ;
 wire \m_blake2.m_hash256.h_flat[130] ;
 wire \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[131] ;
 wire \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[132] ;
 wire \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[133] ;
 wire \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[134] ;
 wire \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[135] ;
 wire \m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[136] ;
 wire \m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[137] ;
 wire \m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[138] ;
 wire \m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[139] ;
 wire \m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[13] ;
 wire \m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2_B1 ;
 wire \m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2_B2 ;
 wire \m_blake2.m_hash256.h_flat[140] ;
 wire \m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[141] ;
 wire \m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[142] ;
 wire \m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[143] ;
 wire \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[144] ;
 wire \m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[145] ;
 wire \m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[146] ;
 wire \m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[147] ;
 wire \m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[148] ;
 wire \m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[149] ;
 wire \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[14] ;
 wire \m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[150] ;
 wire \m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[151] ;
 wire \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[152] ;
 wire \m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[153] ;
 wire \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[154] ;
 wire \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[155] ;
 wire \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[156] ;
 wire \m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[157] ;
 wire \m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[158] ;
 wire \m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[159] ;
 wire \m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[15] ;
 wire \m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[160] ;
 wire \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[161] ;
 wire \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[162] ;
 wire \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[163] ;
 wire \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[164] ;
 wire \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[165] ;
 wire \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[166] ;
 wire \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[167] ;
 wire \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[168] ;
 wire \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[169] ;
 wire \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[16] ;
 wire \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__o22a_2_A2_B1 ;
 wire \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__o22a_2_A2_B2 ;
 wire \m_blake2.m_hash256.h_flat[170] ;
 wire \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[171] ;
 wire \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[172] ;
 wire \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[173] ;
 wire \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[174] ;
 wire \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[175] ;
 wire \m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[176] ;
 wire \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[177] ;
 wire \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[178] ;
 wire \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[179] ;
 wire \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[17] ;
 wire \m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[180] ;
 wire \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[181] ;
 wire \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[182] ;
 wire \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[183] ;
 wire \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[184] ;
 wire \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[185] ;
 wire \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[186] ;
 wire \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[187] ;
 wire \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[188] ;
 wire \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[189] ;
 wire \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[18] ;
 wire \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[190] ;
 wire \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[191] ;
 wire \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[192] ;
 wire \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[193] ;
 wire \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[194] ;
 wire \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[195] ;
 wire \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[196] ;
 wire \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[197] ;
 wire \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[198] ;
 wire \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[199] ;
 wire \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[19] ;
 wire \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_B1 ;
 wire \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_B2 ;
 wire \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[200] ;
 wire \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[201] ;
 wire \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[202] ;
 wire \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[203] ;
 wire \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[204] ;
 wire \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[205] ;
 wire \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[206] ;
 wire \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[207] ;
 wire \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[208] ;
 wire \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[209] ;
 wire \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[20] ;
 wire \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_B1 ;
 wire \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_B2 ;
 wire \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[210] ;
 wire \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[211] ;
 wire \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[212] ;
 wire \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[213] ;
 wire \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[214] ;
 wire \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[215] ;
 wire \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[216] ;
 wire \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[217] ;
 wire \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[218] ;
 wire \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[219] ;
 wire \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[21] ;
 wire \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[220] ;
 wire \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[221] ;
 wire \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[222] ;
 wire \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[223] ;
 wire \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[224] ;
 wire \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[225] ;
 wire \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[226] ;
 wire \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[227] ;
 wire \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[228] ;
 wire \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__a22o_2_A1_B2 ;
 wire \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[229] ;
 wire \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[22] ;
 wire \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[230] ;
 wire \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[231] ;
 wire \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[232] ;
 wire \m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[233] ;
 wire \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[234] ;
 wire \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[235] ;
 wire \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[236] ;
 wire \m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[237] ;
 wire \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[238] ;
 wire \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[239] ;
 wire \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[23] ;
 wire \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[240] ;
 wire \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[241] ;
 wire \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[242] ;
 wire \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[243] ;
 wire \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[244] ;
 wire \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[245] ;
 wire \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[246] ;
 wire \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[247] ;
 wire \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[248] ;
 wire \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__a22o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[249] ;
 wire \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__a22o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[24] ;
 wire \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[250] ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__a22o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__o211a_2_C1_X ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[251] ;
 wire \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__a22o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[252] ;
 wire \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__a22o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[253] ;
 wire \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__a22o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[254] ;
 wire \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__a22o_2_A1_B1 ;
 wire \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[255] ;
 wire \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__a32o_2_B1_A2 ;
 wire \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__a32o_2_B1_A3 ;
 wire \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[25] ;
 wire \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[26] ;
 wire \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[27] ;
 wire \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[28] ;
 wire \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[29] ;
 wire \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[30] ;
 wire \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[31] ;
 wire \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[32] ;
 wire \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[33] ;
 wire \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[34] ;
 wire \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2 ;
 wire \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[35] ;
 wire \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[36] ;
 wire \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[37] ;
 wire \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[38] ;
 wire \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[39] ;
 wire \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[40] ;
 wire \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[41] ;
 wire \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[42] ;
 wire \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[43] ;
 wire \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[44] ;
 wire \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[45] ;
 wire \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[46] ;
 wire \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[47] ;
 wire \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[48] ;
 wire \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[49] ;
 wire \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[50] ;
 wire \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[51] ;
 wire \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[52] ;
 wire \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[53] ;
 wire \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[54] ;
 wire \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[55] ;
 wire \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[56] ;
 wire \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[57] ;
 wire \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[58] ;
 wire \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[59] ;
 wire \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[60] ;
 wire \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[61] ;
 wire \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[62] ;
 wire \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[63] ;
 wire \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[64] ;
 wire \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[65] ;
 wire \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[66] ;
 wire \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[67] ;
 wire \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[68] ;
 wire \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ;
 wire \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[69] ;
 wire \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[70] ;
 wire \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[71] ;
 wire \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[72] ;
 wire \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[73] ;
 wire \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[74] ;
 wire \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[75] ;
 wire \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[76] ;
 wire \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[77] ;
 wire \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[78] ;
 wire \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[79] ;
 wire \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[80] ;
 wire \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ;
 wire \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[81] ;
 wire \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ;
 wire \m_blake2.m_hash256.h_flat[82] ;
 wire \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ;
 wire \m_blake2.m_hash256.h_flat[83] ;
 wire \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[84] ;
 wire \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[85] ;
 wire \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ;
 wire \m_blake2.m_hash256.h_flat[86] ;
 wire \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[87] ;
 wire \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[88] ;
 wire \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[89] ;
 wire \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[8] ;
 wire \m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[90] ;
 wire \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[91] ;
 wire \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[92] ;
 wire \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[93] ;
 wire \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[94] ;
 wire \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[95] ;
 wire \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[96] ;
 wire \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[97] ;
 wire \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[98] ;
 wire \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[99] ;
 wire \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ;
 wire \m_blake2.m_hash256.h_flat[9] ;
 wire \m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ;
 wire \m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.last_block_q ;
 wire \m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a0[0] ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2 ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1 ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[10] ;
 wire \m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[11] ;
 wire \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ;
 wire \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[12] ;
 wire \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[13] ;
 wire \m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[14] ;
 wire \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[15] ;
 wire \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ;
 wire \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2_Y ;
 wire \m_blake2.m_hash256.m_g.a0[16] ;
 wire \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__nor3_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[17] ;
 wire \m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[18] ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a0[19] ;
 wire \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[1] ;
 wire \m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__or3b_2_X_C_N ;
 wire \m_blake2.m_hash256.m_g.a0[20] ;
 wire \m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[21] ;
 wire \m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21bo_2_X_B1_N ;
 wire \m_blake2.m_hash256.m_g.a0[22] ;
 wire \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ;
 wire \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[23] ;
 wire \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[24] ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A3 ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[25] ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_A_N ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1 ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_A1 ;
 wire \m_blake2.m_hash256.m_g.a0[26] ;
 wire \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[27] ;
 wire \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[28] ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ;
 wire \m_blake2.m_hash256.m_g.a0[29] ;
 wire \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[2] ;
 wire \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_A_N ;
 wire \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__or3b_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[30] ;
 wire \m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[31] ;
 wire \m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[3] ;
 wire \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ;
 wire \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[4] ;
 wire \m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[5] ;
 wire \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[6] ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_C_N ;
 wire \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[7] ;
 wire \m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[8] ;
 wire \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.m_g.a0[9] ;
 wire \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.a_q[0] ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[10] ;
 wire \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[11] ;
 wire \m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[12] ;
 wire \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13] ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1_A2 ;
 wire \m_blake2.m_hash256.m_g.a_q[14] ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2 ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[15] ;
 wire \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[16] ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A1 ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A2 ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1 ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[17] ;
 wire \m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[18] ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_A1 ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[19] ;
 wire \m_blake2.m_hash256.m_g.a_q[1] ;
 wire \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[20] ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[21] ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[22] ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A2 ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[23] ;
 wire \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[24] ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[25] ;
 wire \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[26] ;
 wire \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[27] ;
 wire \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.m_g.a_q[28] ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[29] ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_B1 ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X ;
 wire \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[2] ;
 wire \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[30] ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[31] ;
 wire \m_blake2.m_hash256.m_g.a_q[3] ;
 wire \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ba_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[4] ;
 wire \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[5] ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_A2 ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_B ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6] ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_A ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a31o_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[7] ;
 wire \m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[8] ;
 wire \m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9] ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21boi_2_B1_N_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__and3b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[0] ;
 wire \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[10] ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[11] ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1 ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o41a_2_B1_A3 ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12] ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__or4bb_2_C_N_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[13] ;
 wire \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14] ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y_C ;
 wire \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[15] ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16] ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C_X ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__a21o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_B ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[17] ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[18] ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a2111o_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[19] ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[1] ;
 wire \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[20] ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2 ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[21] ;
 wire \m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[22] ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[23] ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_A2 ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[24] ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25] ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A1 ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_A1 ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3 ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B_A ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[26] ;
 wire \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[27] ;
 wire \m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[28] ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_A ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[29] ;
 wire \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[2] ;
 wire \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[30] ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1 ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3 ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2 ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[31] ;
 wire \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ;
 wire \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[3] ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[4] ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_B ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5] ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[6] ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_A2 ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[7] ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[8] ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.b_q[9] ;
 wire \m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[0] ;
 wire \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[10] ;
 wire \m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[11] ;
 wire \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[12] ;
 wire \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[13] ;
 wire \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[14] ;
 wire \m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[15] ;
 wire \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_A4 ;
 wire \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__o211a_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[16] ;
 wire \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_B ;
 wire \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[17] ;
 wire \m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[18] ;
 wire \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[19] ;
 wire \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B2 ;
 wire \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__o211a_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[1] ;
 wire \m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[20] ;
 wire \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[21] ;
 wire \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[22] ;
 wire \m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[23] ;
 wire \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ;
 wire \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[24] ;
 wire \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[25] ;
 wire \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[26] ;
 wire \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[27] ;
 wire \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ;
 wire \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X ;
 wire \m_blake2.m_hash256.m_g.c_q[28] ;
 wire \m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[29] ;
 wire \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[2] ;
 wire \m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[30] ;
 wire \m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[31] ;
 wire \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_B ;
 wire \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[3] ;
 wire \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B2 ;
 wire \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__o211a_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[4] ;
 wire \m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[5] ;
 wire \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[6] ;
 wire \m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[7] ;
 wire \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_A2 ;
 wire \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_B1 ;
 wire \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_X ;
 wire \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__o21bai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.c_q[8] ;
 wire \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[9] ;
 wire \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.d_q[0] ;
 wire \m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[10] ;
 wire \m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[11] ;
 wire \m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[12] ;
 wire \m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[13] ;
 wire \m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[14] ;
 wire \m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[15] ;
 wire \m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.d_q[16] ;
 wire \m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[17] ;
 wire \m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[18] ;
 wire \m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[19] ;
 wire \m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[1] ;
 wire \m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[20] ;
 wire \m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[21] ;
 wire \m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[22] ;
 wire \m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[23] ;
 wire \m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[24] ;
 wire \m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[25] ;
 wire \m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[26] ;
 wire \m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[27] ;
 wire \m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[28] ;
 wire \m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[29] ;
 wire \m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[2] ;
 wire \m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[30] ;
 wire \m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[31] ;
 wire \m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[3] ;
 wire \m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[4] ;
 wire \m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[5] ;
 wire \m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[6] ;
 wire \m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[7] ;
 wire \m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[8] ;
 wire \m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.d_q[9] ;
 wire \m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[0] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[10] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[11] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[12] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[13] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[14] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[15] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[16] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[17] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[18] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[19] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[1] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[20] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[21] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[22] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[23] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2_B1 ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[25] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[26] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[27] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[28] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[29] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[2] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[30] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[31] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[31]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[3] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[4] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[5] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[6] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[8] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[9] ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.m_matrix[0][0] ;
 wire \m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_blake2.m_hash256.m_matrix[0][10] ;
 wire \m_blake2.m_hash256.m_matrix[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][11] ;
 wire \m_blake2.m_hash256.m_matrix[0][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][12] ;
 wire \m_blake2.m_hash256.m_matrix[0][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][13] ;
 wire \m_blake2.m_hash256.m_matrix[0][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][14] ;
 wire \m_blake2.m_hash256.m_matrix[0][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][15] ;
 wire \m_blake2.m_hash256.m_matrix[0][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][16] ;
 wire \m_blake2.m_hash256.m_matrix[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][17] ;
 wire \m_blake2.m_hash256.m_matrix[0][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][18] ;
 wire \m_blake2.m_hash256.m_matrix[0][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][19] ;
 wire \m_blake2.m_hash256.m_matrix[0][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][1] ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1 ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2 ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3 ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X ;
 wire \m_blake2.m_hash256.m_matrix[0][20] ;
 wire \m_blake2.m_hash256.m_matrix[0][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][21] ;
 wire \m_blake2.m_hash256.m_matrix[0][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][22] ;
 wire \m_blake2.m_hash256.m_matrix[0][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][23] ;
 wire \m_blake2.m_hash256.m_matrix[0][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][24] ;
 wire \m_blake2.m_hash256.m_matrix[0][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][25] ;
 wire \m_blake2.m_hash256.m_matrix[0][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][26] ;
 wire \m_blake2.m_hash256.m_matrix[0][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][27] ;
 wire \m_blake2.m_hash256.m_matrix[0][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][28] ;
 wire \m_blake2.m_hash256.m_matrix[0][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][29] ;
 wire \m_blake2.m_hash256.m_matrix[0][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][2] ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1 ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2 ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3 ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X ;
 wire \m_blake2.m_hash256.m_matrix[0][30] ;
 wire \m_blake2.m_hash256.m_matrix[0][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][31] ;
 wire \m_blake2.m_hash256.m_matrix[0][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][3] ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2 ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X ;
 wire \m_blake2.m_hash256.m_matrix[0][4] ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_matrix[0][5] ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2 ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_matrix[0][6] ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2 ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X ;
 wire \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.m_matrix[0][7] ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y ;
 wire \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_X ;
 wire \m_blake2.m_hash256.m_matrix[0][8] ;
 wire \m_blake2.m_hash256.m_matrix[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[0][9] ;
 wire \m_blake2.m_hash256.m_matrix[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][0] ;
 wire \m_blake2.m_hash256.m_matrix[10][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][10] ;
 wire \m_blake2.m_hash256.m_matrix[10][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][11] ;
 wire \m_blake2.m_hash256.m_matrix[10][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][12] ;
 wire \m_blake2.m_hash256.m_matrix[10][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][13] ;
 wire \m_blake2.m_hash256.m_matrix[10][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][14] ;
 wire \m_blake2.m_hash256.m_matrix[10][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][15] ;
 wire \m_blake2.m_hash256.m_matrix[10][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][16] ;
 wire \m_blake2.m_hash256.m_matrix[10][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][17] ;
 wire \m_blake2.m_hash256.m_matrix[10][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][18] ;
 wire \m_blake2.m_hash256.m_matrix[10][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][19] ;
 wire \m_blake2.m_hash256.m_matrix[10][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][1] ;
 wire \m_blake2.m_hash256.m_matrix[10][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][20] ;
 wire \m_blake2.m_hash256.m_matrix[10][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][21] ;
 wire \m_blake2.m_hash256.m_matrix[10][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][22] ;
 wire \m_blake2.m_hash256.m_matrix[10][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][23] ;
 wire \m_blake2.m_hash256.m_matrix[10][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][24] ;
 wire \m_blake2.m_hash256.m_matrix[10][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][25] ;
 wire \m_blake2.m_hash256.m_matrix[10][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][26] ;
 wire \m_blake2.m_hash256.m_matrix[10][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][27] ;
 wire \m_blake2.m_hash256.m_matrix[10][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][28] ;
 wire \m_blake2.m_hash256.m_matrix[10][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][29] ;
 wire \m_blake2.m_hash256.m_matrix[10][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][2] ;
 wire \m_blake2.m_hash256.m_matrix[10][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][30] ;
 wire \m_blake2.m_hash256.m_matrix[10][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][31] ;
 wire \m_blake2.m_hash256.m_matrix[10][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][3] ;
 wire \m_blake2.m_hash256.m_matrix[10][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][4] ;
 wire \m_blake2.m_hash256.m_matrix[10][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][5] ;
 wire \m_blake2.m_hash256.m_matrix[10][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][6] ;
 wire \m_blake2.m_hash256.m_matrix[10][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][7] ;
 wire \m_blake2.m_hash256.m_matrix[10][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][8] ;
 wire \m_blake2.m_hash256.m_matrix[10][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[10][9] ;
 wire \m_blake2.m_hash256.m_matrix[10][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][0] ;
 wire \m_blake2.m_hash256.m_matrix[11][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][10] ;
 wire \m_blake2.m_hash256.m_matrix[11][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][11] ;
 wire \m_blake2.m_hash256.m_matrix[11][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][12] ;
 wire \m_blake2.m_hash256.m_matrix[11][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][13] ;
 wire \m_blake2.m_hash256.m_matrix[11][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][14] ;
 wire \m_blake2.m_hash256.m_matrix[11][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][15] ;
 wire \m_blake2.m_hash256.m_matrix[11][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][16] ;
 wire \m_blake2.m_hash256.m_matrix[11][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][17] ;
 wire \m_blake2.m_hash256.m_matrix[11][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][18] ;
 wire \m_blake2.m_hash256.m_matrix[11][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][19] ;
 wire \m_blake2.m_hash256.m_matrix[11][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][1] ;
 wire \m_blake2.m_hash256.m_matrix[11][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][20] ;
 wire \m_blake2.m_hash256.m_matrix[11][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][21] ;
 wire \m_blake2.m_hash256.m_matrix[11][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][22] ;
 wire \m_blake2.m_hash256.m_matrix[11][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][23] ;
 wire \m_blake2.m_hash256.m_matrix[11][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][24] ;
 wire \m_blake2.m_hash256.m_matrix[11][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][25] ;
 wire \m_blake2.m_hash256.m_matrix[11][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][26] ;
 wire \m_blake2.m_hash256.m_matrix[11][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][27] ;
 wire \m_blake2.m_hash256.m_matrix[11][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][28] ;
 wire \m_blake2.m_hash256.m_matrix[11][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][29] ;
 wire \m_blake2.m_hash256.m_matrix[11][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][2] ;
 wire \m_blake2.m_hash256.m_matrix[11][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][30] ;
 wire \m_blake2.m_hash256.m_matrix[11][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][31] ;
 wire \m_blake2.m_hash256.m_matrix[11][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][3] ;
 wire \m_blake2.m_hash256.m_matrix[11][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][4] ;
 wire \m_blake2.m_hash256.m_matrix[11][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][5] ;
 wire \m_blake2.m_hash256.m_matrix[11][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][6] ;
 wire \m_blake2.m_hash256.m_matrix[11][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][7] ;
 wire \m_blake2.m_hash256.m_matrix[11][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][8] ;
 wire \m_blake2.m_hash256.m_matrix[11][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[11][9] ;
 wire \m_blake2.m_hash256.m_matrix[11][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][0] ;
 wire \m_blake2.m_hash256.m_matrix[12][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][10] ;
 wire \m_blake2.m_hash256.m_matrix[12][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][11] ;
 wire \m_blake2.m_hash256.m_matrix[12][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][12] ;
 wire \m_blake2.m_hash256.m_matrix[12][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][13] ;
 wire \m_blake2.m_hash256.m_matrix[12][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][14] ;
 wire \m_blake2.m_hash256.m_matrix[12][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][15] ;
 wire \m_blake2.m_hash256.m_matrix[12][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][16] ;
 wire \m_blake2.m_hash256.m_matrix[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][17] ;
 wire \m_blake2.m_hash256.m_matrix[12][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][18] ;
 wire \m_blake2.m_hash256.m_matrix[12][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][19] ;
 wire \m_blake2.m_hash256.m_matrix[12][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][1] ;
 wire \m_blake2.m_hash256.m_matrix[12][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][20] ;
 wire \m_blake2.m_hash256.m_matrix[12][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][21] ;
 wire \m_blake2.m_hash256.m_matrix[12][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][22] ;
 wire \m_blake2.m_hash256.m_matrix[12][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][23] ;
 wire \m_blake2.m_hash256.m_matrix[12][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][24] ;
 wire \m_blake2.m_hash256.m_matrix[12][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][25] ;
 wire \m_blake2.m_hash256.m_matrix[12][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][26] ;
 wire \m_blake2.m_hash256.m_matrix[12][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][27] ;
 wire \m_blake2.m_hash256.m_matrix[12][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][28] ;
 wire \m_blake2.m_hash256.m_matrix[12][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][29] ;
 wire \m_blake2.m_hash256.m_matrix[12][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][2] ;
 wire \m_blake2.m_hash256.m_matrix[12][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][30] ;
 wire \m_blake2.m_hash256.m_matrix[12][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][31] ;
 wire \m_blake2.m_hash256.m_matrix[12][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][3] ;
 wire \m_blake2.m_hash256.m_matrix[12][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][4] ;
 wire \m_blake2.m_hash256.m_matrix[12][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][5] ;
 wire \m_blake2.m_hash256.m_matrix[12][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][6] ;
 wire \m_blake2.m_hash256.m_matrix[12][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][7] ;
 wire \m_blake2.m_hash256.m_matrix[12][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][8] ;
 wire \m_blake2.m_hash256.m_matrix[12][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[12][9] ;
 wire \m_blake2.m_hash256.m_matrix[12][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][0] ;
 wire \m_blake2.m_hash256.m_matrix[13][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][10] ;
 wire \m_blake2.m_hash256.m_matrix[13][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][11] ;
 wire \m_blake2.m_hash256.m_matrix[13][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][12] ;
 wire \m_blake2.m_hash256.m_matrix[13][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][13] ;
 wire \m_blake2.m_hash256.m_matrix[13][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][14] ;
 wire \m_blake2.m_hash256.m_matrix[13][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][15] ;
 wire \m_blake2.m_hash256.m_matrix[13][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][16] ;
 wire \m_blake2.m_hash256.m_matrix[13][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][17] ;
 wire \m_blake2.m_hash256.m_matrix[13][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][18] ;
 wire \m_blake2.m_hash256.m_matrix[13][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][19] ;
 wire \m_blake2.m_hash256.m_matrix[13][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][1] ;
 wire \m_blake2.m_hash256.m_matrix[13][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][20] ;
 wire \m_blake2.m_hash256.m_matrix[13][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][21] ;
 wire \m_blake2.m_hash256.m_matrix[13][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][22] ;
 wire \m_blake2.m_hash256.m_matrix[13][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][23] ;
 wire \m_blake2.m_hash256.m_matrix[13][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][24] ;
 wire \m_blake2.m_hash256.m_matrix[13][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][25] ;
 wire \m_blake2.m_hash256.m_matrix[13][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][26] ;
 wire \m_blake2.m_hash256.m_matrix[13][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][27] ;
 wire \m_blake2.m_hash256.m_matrix[13][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][28] ;
 wire \m_blake2.m_hash256.m_matrix[13][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][29] ;
 wire \m_blake2.m_hash256.m_matrix[13][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][2] ;
 wire \m_blake2.m_hash256.m_matrix[13][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][30] ;
 wire \m_blake2.m_hash256.m_matrix[13][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][31] ;
 wire \m_blake2.m_hash256.m_matrix[13][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][3] ;
 wire \m_blake2.m_hash256.m_matrix[13][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][4] ;
 wire \m_blake2.m_hash256.m_matrix[13][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][5] ;
 wire \m_blake2.m_hash256.m_matrix[13][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][6] ;
 wire \m_blake2.m_hash256.m_matrix[13][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][7] ;
 wire \m_blake2.m_hash256.m_matrix[13][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][8] ;
 wire \m_blake2.m_hash256.m_matrix[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[13][9] ;
 wire \m_blake2.m_hash256.m_matrix[13][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][0] ;
 wire \m_blake2.m_hash256.m_matrix[14][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][10] ;
 wire \m_blake2.m_hash256.m_matrix[14][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][11] ;
 wire \m_blake2.m_hash256.m_matrix[14][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][12] ;
 wire \m_blake2.m_hash256.m_matrix[14][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][13] ;
 wire \m_blake2.m_hash256.m_matrix[14][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][14] ;
 wire \m_blake2.m_hash256.m_matrix[14][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][15] ;
 wire \m_blake2.m_hash256.m_matrix[14][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][16] ;
 wire \m_blake2.m_hash256.m_matrix[14][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][17] ;
 wire \m_blake2.m_hash256.m_matrix[14][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][18] ;
 wire \m_blake2.m_hash256.m_matrix[14][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][19] ;
 wire \m_blake2.m_hash256.m_matrix[14][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][1] ;
 wire \m_blake2.m_hash256.m_matrix[14][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][20] ;
 wire \m_blake2.m_hash256.m_matrix[14][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][21] ;
 wire \m_blake2.m_hash256.m_matrix[14][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][22] ;
 wire \m_blake2.m_hash256.m_matrix[14][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][23] ;
 wire \m_blake2.m_hash256.m_matrix[14][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][24] ;
 wire \m_blake2.m_hash256.m_matrix[14][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][25] ;
 wire \m_blake2.m_hash256.m_matrix[14][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][26] ;
 wire \m_blake2.m_hash256.m_matrix[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][27] ;
 wire \m_blake2.m_hash256.m_matrix[14][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][28] ;
 wire \m_blake2.m_hash256.m_matrix[14][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][29] ;
 wire \m_blake2.m_hash256.m_matrix[14][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][2] ;
 wire \m_blake2.m_hash256.m_matrix[14][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][30] ;
 wire \m_blake2.m_hash256.m_matrix[14][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][31] ;
 wire \m_blake2.m_hash256.m_matrix[14][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][3] ;
 wire \m_blake2.m_hash256.m_matrix[14][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][4] ;
 wire \m_blake2.m_hash256.m_matrix[14][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][5] ;
 wire \m_blake2.m_hash256.m_matrix[14][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][6] ;
 wire \m_blake2.m_hash256.m_matrix[14][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][7] ;
 wire \m_blake2.m_hash256.m_matrix[14][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][8] ;
 wire \m_blake2.m_hash256.m_matrix[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[14][9] ;
 wire \m_blake2.m_hash256.m_matrix[14][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][0] ;
 wire \m_blake2.m_hash256.m_matrix[15][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][10] ;
 wire \m_blake2.m_hash256.m_matrix[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][11] ;
 wire \m_blake2.m_hash256.m_matrix[15][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][12] ;
 wire \m_blake2.m_hash256.m_matrix[15][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][13] ;
 wire \m_blake2.m_hash256.m_matrix[15][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][14] ;
 wire \m_blake2.m_hash256.m_matrix[15][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][15] ;
 wire \m_blake2.m_hash256.m_matrix[15][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][16] ;
 wire \m_blake2.m_hash256.m_matrix[15][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][17] ;
 wire \m_blake2.m_hash256.m_matrix[15][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][18] ;
 wire \m_blake2.m_hash256.m_matrix[15][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][19] ;
 wire \m_blake2.m_hash256.m_matrix[15][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][1] ;
 wire \m_blake2.m_hash256.m_matrix[15][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][20] ;
 wire \m_blake2.m_hash256.m_matrix[15][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][21] ;
 wire \m_blake2.m_hash256.m_matrix[15][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][22] ;
 wire \m_blake2.m_hash256.m_matrix[15][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][23] ;
 wire \m_blake2.m_hash256.m_matrix[15][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][24] ;
 wire \m_blake2.m_hash256.m_matrix[15][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][25] ;
 wire \m_blake2.m_hash256.m_matrix[15][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][26] ;
 wire \m_blake2.m_hash256.m_matrix[15][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][27] ;
 wire \m_blake2.m_hash256.m_matrix[15][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][28] ;
 wire \m_blake2.m_hash256.m_matrix[15][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][29] ;
 wire \m_blake2.m_hash256.m_matrix[15][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][2] ;
 wire \m_blake2.m_hash256.m_matrix[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][30] ;
 wire \m_blake2.m_hash256.m_matrix[15][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][31] ;
 wire \m_blake2.m_hash256.m_matrix[15][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][3] ;
 wire \m_blake2.m_hash256.m_matrix[15][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][4] ;
 wire \m_blake2.m_hash256.m_matrix[15][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][5] ;
 wire \m_blake2.m_hash256.m_matrix[15][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][6] ;
 wire \m_blake2.m_hash256.m_matrix[15][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][7] ;
 wire \m_blake2.m_hash256.m_matrix[15][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][8] ;
 wire \m_blake2.m_hash256.m_matrix[15][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[15][9] ;
 wire \m_blake2.m_hash256.m_matrix[15][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][0] ;
 wire \m_blake2.m_hash256.m_matrix[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][10] ;
 wire \m_blake2.m_hash256.m_matrix[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][11] ;
 wire \m_blake2.m_hash256.m_matrix[1][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][12] ;
 wire \m_blake2.m_hash256.m_matrix[1][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][13] ;
 wire \m_blake2.m_hash256.m_matrix[1][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][14] ;
 wire \m_blake2.m_hash256.m_matrix[1][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][15] ;
 wire \m_blake2.m_hash256.m_matrix[1][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][16] ;
 wire \m_blake2.m_hash256.m_matrix[1][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][17] ;
 wire \m_blake2.m_hash256.m_matrix[1][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][18] ;
 wire \m_blake2.m_hash256.m_matrix[1][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][19] ;
 wire \m_blake2.m_hash256.m_matrix[1][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][1] ;
 wire \m_blake2.m_hash256.m_matrix[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][20] ;
 wire \m_blake2.m_hash256.m_matrix[1][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][21] ;
 wire \m_blake2.m_hash256.m_matrix[1][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][22] ;
 wire \m_blake2.m_hash256.m_matrix[1][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][23] ;
 wire \m_blake2.m_hash256.m_matrix[1][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][24] ;
 wire \m_blake2.m_hash256.m_matrix[1][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][25] ;
 wire \m_blake2.m_hash256.m_matrix[1][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][26] ;
 wire \m_blake2.m_hash256.m_matrix[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][27] ;
 wire \m_blake2.m_hash256.m_matrix[1][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][28] ;
 wire \m_blake2.m_hash256.m_matrix[1][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][29] ;
 wire \m_blake2.m_hash256.m_matrix[1][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][2] ;
 wire \m_blake2.m_hash256.m_matrix[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][30] ;
 wire \m_blake2.m_hash256.m_matrix[1][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][31] ;
 wire \m_blake2.m_hash256.m_matrix[1][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][3] ;
 wire \m_blake2.m_hash256.m_matrix[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][4] ;
 wire \m_blake2.m_hash256.m_matrix[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][5] ;
 wire \m_blake2.m_hash256.m_matrix[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][6] ;
 wire \m_blake2.m_hash256.m_matrix[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][7] ;
 wire \m_blake2.m_hash256.m_matrix[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][8] ;
 wire \m_blake2.m_hash256.m_matrix[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[1][9] ;
 wire \m_blake2.m_hash256.m_matrix[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][0] ;
 wire \m_blake2.m_hash256.m_matrix[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][10] ;
 wire \m_blake2.m_hash256.m_matrix[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][11] ;
 wire \m_blake2.m_hash256.m_matrix[2][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][12] ;
 wire \m_blake2.m_hash256.m_matrix[2][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][13] ;
 wire \m_blake2.m_hash256.m_matrix[2][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][14] ;
 wire \m_blake2.m_hash256.m_matrix[2][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][15] ;
 wire \m_blake2.m_hash256.m_matrix[2][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][16] ;
 wire \m_blake2.m_hash256.m_matrix[2][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][17] ;
 wire \m_blake2.m_hash256.m_matrix[2][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][18] ;
 wire \m_blake2.m_hash256.m_matrix[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][19] ;
 wire \m_blake2.m_hash256.m_matrix[2][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][1] ;
 wire \m_blake2.m_hash256.m_matrix[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][20] ;
 wire \m_blake2.m_hash256.m_matrix[2][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][21] ;
 wire \m_blake2.m_hash256.m_matrix[2][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][22] ;
 wire \m_blake2.m_hash256.m_matrix[2][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][23] ;
 wire \m_blake2.m_hash256.m_matrix[2][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][24] ;
 wire \m_blake2.m_hash256.m_matrix[2][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][25] ;
 wire \m_blake2.m_hash256.m_matrix[2][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][26] ;
 wire \m_blake2.m_hash256.m_matrix[2][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][27] ;
 wire \m_blake2.m_hash256.m_matrix[2][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][28] ;
 wire \m_blake2.m_hash256.m_matrix[2][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][29] ;
 wire \m_blake2.m_hash256.m_matrix[2][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][2] ;
 wire \m_blake2.m_hash256.m_matrix[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][30] ;
 wire \m_blake2.m_hash256.m_matrix[2][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][31] ;
 wire \m_blake2.m_hash256.m_matrix[2][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][3] ;
 wire \m_blake2.m_hash256.m_matrix[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][4] ;
 wire \m_blake2.m_hash256.m_matrix[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][5] ;
 wire \m_blake2.m_hash256.m_matrix[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][6] ;
 wire \m_blake2.m_hash256.m_matrix[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][7] ;
 wire \m_blake2.m_hash256.m_matrix[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][8] ;
 wire \m_blake2.m_hash256.m_matrix[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[2][9] ;
 wire \m_blake2.m_hash256.m_matrix[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][0] ;
 wire \m_blake2.m_hash256.m_matrix[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][10] ;
 wire \m_blake2.m_hash256.m_matrix[3][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][11] ;
 wire \m_blake2.m_hash256.m_matrix[3][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][12] ;
 wire \m_blake2.m_hash256.m_matrix[3][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][13] ;
 wire \m_blake2.m_hash256.m_matrix[3][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][14] ;
 wire \m_blake2.m_hash256.m_matrix[3][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][15] ;
 wire \m_blake2.m_hash256.m_matrix[3][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][16] ;
 wire \m_blake2.m_hash256.m_matrix[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][17] ;
 wire \m_blake2.m_hash256.m_matrix[3][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][18] ;
 wire \m_blake2.m_hash256.m_matrix[3][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][19] ;
 wire \m_blake2.m_hash256.m_matrix[3][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][1] ;
 wire \m_blake2.m_hash256.m_matrix[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][20] ;
 wire \m_blake2.m_hash256.m_matrix[3][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][21] ;
 wire \m_blake2.m_hash256.m_matrix[3][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][22] ;
 wire \m_blake2.m_hash256.m_matrix[3][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][23] ;
 wire \m_blake2.m_hash256.m_matrix[3][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][24] ;
 wire \m_blake2.m_hash256.m_matrix[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][25] ;
 wire \m_blake2.m_hash256.m_matrix[3][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][26] ;
 wire \m_blake2.m_hash256.m_matrix[3][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][27] ;
 wire \m_blake2.m_hash256.m_matrix[3][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][28] ;
 wire \m_blake2.m_hash256.m_matrix[3][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][29] ;
 wire \m_blake2.m_hash256.m_matrix[3][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][2] ;
 wire \m_blake2.m_hash256.m_matrix[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][30] ;
 wire \m_blake2.m_hash256.m_matrix[3][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][31] ;
 wire \m_blake2.m_hash256.m_matrix[3][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][3] ;
 wire \m_blake2.m_hash256.m_matrix[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][4] ;
 wire \m_blake2.m_hash256.m_matrix[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][5] ;
 wire \m_blake2.m_hash256.m_matrix[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][6] ;
 wire \m_blake2.m_hash256.m_matrix[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][7] ;
 wire \m_blake2.m_hash256.m_matrix[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][8] ;
 wire \m_blake2.m_hash256.m_matrix[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[3][9] ;
 wire \m_blake2.m_hash256.m_matrix[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][0] ;
 wire \m_blake2.m_hash256.m_matrix[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][10] ;
 wire \m_blake2.m_hash256.m_matrix[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][11] ;
 wire \m_blake2.m_hash256.m_matrix[4][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][12] ;
 wire \m_blake2.m_hash256.m_matrix[4][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][13] ;
 wire \m_blake2.m_hash256.m_matrix[4][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][14] ;
 wire \m_blake2.m_hash256.m_matrix[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][15] ;
 wire \m_blake2.m_hash256.m_matrix[4][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][16] ;
 wire \m_blake2.m_hash256.m_matrix[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][17] ;
 wire \m_blake2.m_hash256.m_matrix[4][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][18] ;
 wire \m_blake2.m_hash256.m_matrix[4][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][19] ;
 wire \m_blake2.m_hash256.m_matrix[4][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][1] ;
 wire \m_blake2.m_hash256.m_matrix[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][20] ;
 wire \m_blake2.m_hash256.m_matrix[4][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][21] ;
 wire \m_blake2.m_hash256.m_matrix[4][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][22] ;
 wire \m_blake2.m_hash256.m_matrix[4][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][23] ;
 wire \m_blake2.m_hash256.m_matrix[4][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][24] ;
 wire \m_blake2.m_hash256.m_matrix[4][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][25] ;
 wire \m_blake2.m_hash256.m_matrix[4][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][26] ;
 wire \m_blake2.m_hash256.m_matrix[4][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][27] ;
 wire \m_blake2.m_hash256.m_matrix[4][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][28] ;
 wire \m_blake2.m_hash256.m_matrix[4][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][29] ;
 wire \m_blake2.m_hash256.m_matrix[4][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][2] ;
 wire \m_blake2.m_hash256.m_matrix[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][30] ;
 wire \m_blake2.m_hash256.m_matrix[4][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][31] ;
 wire \m_blake2.m_hash256.m_matrix[4][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][3] ;
 wire \m_blake2.m_hash256.m_matrix[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][4] ;
 wire \m_blake2.m_hash256.m_matrix[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][5] ;
 wire \m_blake2.m_hash256.m_matrix[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][6] ;
 wire \m_blake2.m_hash256.m_matrix[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][7] ;
 wire \m_blake2.m_hash256.m_matrix[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][8] ;
 wire \m_blake2.m_hash256.m_matrix[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[4][9] ;
 wire \m_blake2.m_hash256.m_matrix[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][0] ;
 wire \m_blake2.m_hash256.m_matrix[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][10] ;
 wire \m_blake2.m_hash256.m_matrix[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][11] ;
 wire \m_blake2.m_hash256.m_matrix[5][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][12] ;
 wire \m_blake2.m_hash256.m_matrix[5][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][13] ;
 wire \m_blake2.m_hash256.m_matrix[5][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][14] ;
 wire \m_blake2.m_hash256.m_matrix[5][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][15] ;
 wire \m_blake2.m_hash256.m_matrix[5][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][16] ;
 wire \m_blake2.m_hash256.m_matrix[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][17] ;
 wire \m_blake2.m_hash256.m_matrix[5][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][18] ;
 wire \m_blake2.m_hash256.m_matrix[5][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][19] ;
 wire \m_blake2.m_hash256.m_matrix[5][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][1] ;
 wire \m_blake2.m_hash256.m_matrix[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][20] ;
 wire \m_blake2.m_hash256.m_matrix[5][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][21] ;
 wire \m_blake2.m_hash256.m_matrix[5][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][22] ;
 wire \m_blake2.m_hash256.m_matrix[5][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][23] ;
 wire \m_blake2.m_hash256.m_matrix[5][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][24] ;
 wire \m_blake2.m_hash256.m_matrix[5][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][25] ;
 wire \m_blake2.m_hash256.m_matrix[5][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][26] ;
 wire \m_blake2.m_hash256.m_matrix[5][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][27] ;
 wire \m_blake2.m_hash256.m_matrix[5][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][28] ;
 wire \m_blake2.m_hash256.m_matrix[5][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][29] ;
 wire \m_blake2.m_hash256.m_matrix[5][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][2] ;
 wire \m_blake2.m_hash256.m_matrix[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][30] ;
 wire \m_blake2.m_hash256.m_matrix[5][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][31] ;
 wire \m_blake2.m_hash256.m_matrix[5][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][3] ;
 wire \m_blake2.m_hash256.m_matrix[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][4] ;
 wire \m_blake2.m_hash256.m_matrix[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][5] ;
 wire \m_blake2.m_hash256.m_matrix[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][6] ;
 wire \m_blake2.m_hash256.m_matrix[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][7] ;
 wire \m_blake2.m_hash256.m_matrix[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][8] ;
 wire \m_blake2.m_hash256.m_matrix[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[5][9] ;
 wire \m_blake2.m_hash256.m_matrix[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][0] ;
 wire \m_blake2.m_hash256.m_matrix[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][10] ;
 wire \m_blake2.m_hash256.m_matrix[6][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][11] ;
 wire \m_blake2.m_hash256.m_matrix[6][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][12] ;
 wire \m_blake2.m_hash256.m_matrix[6][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][13] ;
 wire \m_blake2.m_hash256.m_matrix[6][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][14] ;
 wire \m_blake2.m_hash256.m_matrix[6][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][15] ;
 wire \m_blake2.m_hash256.m_matrix[6][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][16] ;
 wire \m_blake2.m_hash256.m_matrix[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][17] ;
 wire \m_blake2.m_hash256.m_matrix[6][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][18] ;
 wire \m_blake2.m_hash256.m_matrix[6][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][19] ;
 wire \m_blake2.m_hash256.m_matrix[6][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][1] ;
 wire \m_blake2.m_hash256.m_matrix[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][20] ;
 wire \m_blake2.m_hash256.m_matrix[6][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][21] ;
 wire \m_blake2.m_hash256.m_matrix[6][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][22] ;
 wire \m_blake2.m_hash256.m_matrix[6][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][23] ;
 wire \m_blake2.m_hash256.m_matrix[6][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][24] ;
 wire \m_blake2.m_hash256.m_matrix[6][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][25] ;
 wire \m_blake2.m_hash256.m_matrix[6][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][26] ;
 wire \m_blake2.m_hash256.m_matrix[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][27] ;
 wire \m_blake2.m_hash256.m_matrix[6][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][28] ;
 wire \m_blake2.m_hash256.m_matrix[6][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][29] ;
 wire \m_blake2.m_hash256.m_matrix[6][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][2] ;
 wire \m_blake2.m_hash256.m_matrix[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][30] ;
 wire \m_blake2.m_hash256.m_matrix[6][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][31] ;
 wire \m_blake2.m_hash256.m_matrix[6][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][3] ;
 wire \m_blake2.m_hash256.m_matrix[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][4] ;
 wire \m_blake2.m_hash256.m_matrix[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][5] ;
 wire \m_blake2.m_hash256.m_matrix[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][6] ;
 wire \m_blake2.m_hash256.m_matrix[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][7] ;
 wire \m_blake2.m_hash256.m_matrix[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][8] ;
 wire \m_blake2.m_hash256.m_matrix[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[6][9] ;
 wire \m_blake2.m_hash256.m_matrix[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][0] ;
 wire \m_blake2.m_hash256.m_matrix[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][10] ;
 wire \m_blake2.m_hash256.m_matrix[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][11] ;
 wire \m_blake2.m_hash256.m_matrix[7][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][12] ;
 wire \m_blake2.m_hash256.m_matrix[7][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][13] ;
 wire \m_blake2.m_hash256.m_matrix[7][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][14] ;
 wire \m_blake2.m_hash256.m_matrix[7][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][15] ;
 wire \m_blake2.m_hash256.m_matrix[7][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][16] ;
 wire \m_blake2.m_hash256.m_matrix[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][17] ;
 wire \m_blake2.m_hash256.m_matrix[7][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][18] ;
 wire \m_blake2.m_hash256.m_matrix[7][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][19] ;
 wire \m_blake2.m_hash256.m_matrix[7][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][1] ;
 wire \m_blake2.m_hash256.m_matrix[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][20] ;
 wire \m_blake2.m_hash256.m_matrix[7][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][21] ;
 wire \m_blake2.m_hash256.m_matrix[7][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][22] ;
 wire \m_blake2.m_hash256.m_matrix[7][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][23] ;
 wire \m_blake2.m_hash256.m_matrix[7][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][24] ;
 wire \m_blake2.m_hash256.m_matrix[7][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][25] ;
 wire \m_blake2.m_hash256.m_matrix[7][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][26] ;
 wire \m_blake2.m_hash256.m_matrix[7][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][27] ;
 wire \m_blake2.m_hash256.m_matrix[7][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][28] ;
 wire \m_blake2.m_hash256.m_matrix[7][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][29] ;
 wire \m_blake2.m_hash256.m_matrix[7][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][2] ;
 wire \m_blake2.m_hash256.m_matrix[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][30] ;
 wire \m_blake2.m_hash256.m_matrix[7][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][31] ;
 wire \m_blake2.m_hash256.m_matrix[7][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][3] ;
 wire \m_blake2.m_hash256.m_matrix[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][4] ;
 wire \m_blake2.m_hash256.m_matrix[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][5] ;
 wire \m_blake2.m_hash256.m_matrix[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][6] ;
 wire \m_blake2.m_hash256.m_matrix[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][7] ;
 wire \m_blake2.m_hash256.m_matrix[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][8] ;
 wire \m_blake2.m_hash256.m_matrix[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[7][9] ;
 wire \m_blake2.m_hash256.m_matrix[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][0] ;
 wire \m_blake2.m_hash256.m_matrix[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][10] ;
 wire \m_blake2.m_hash256.m_matrix[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][11] ;
 wire \m_blake2.m_hash256.m_matrix[8][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][12] ;
 wire \m_blake2.m_hash256.m_matrix[8][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][13] ;
 wire \m_blake2.m_hash256.m_matrix[8][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][14] ;
 wire \m_blake2.m_hash256.m_matrix[8][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][15] ;
 wire \m_blake2.m_hash256.m_matrix[8][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][16] ;
 wire \m_blake2.m_hash256.m_matrix[8][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][17] ;
 wire \m_blake2.m_hash256.m_matrix[8][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][18] ;
 wire \m_blake2.m_hash256.m_matrix[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][19] ;
 wire \m_blake2.m_hash256.m_matrix[8][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][1] ;
 wire \m_blake2.m_hash256.m_matrix[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][20] ;
 wire \m_blake2.m_hash256.m_matrix[8][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][21] ;
 wire \m_blake2.m_hash256.m_matrix[8][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][22] ;
 wire \m_blake2.m_hash256.m_matrix[8][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][23] ;
 wire \m_blake2.m_hash256.m_matrix[8][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][24] ;
 wire \m_blake2.m_hash256.m_matrix[8][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][25] ;
 wire \m_blake2.m_hash256.m_matrix[8][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][26] ;
 wire \m_blake2.m_hash256.m_matrix[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][27] ;
 wire \m_blake2.m_hash256.m_matrix[8][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][28] ;
 wire \m_blake2.m_hash256.m_matrix[8][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][29] ;
 wire \m_blake2.m_hash256.m_matrix[8][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][2] ;
 wire \m_blake2.m_hash256.m_matrix[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][30] ;
 wire \m_blake2.m_hash256.m_matrix[8][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][31] ;
 wire \m_blake2.m_hash256.m_matrix[8][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][3] ;
 wire \m_blake2.m_hash256.m_matrix[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][4] ;
 wire \m_blake2.m_hash256.m_matrix[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][5] ;
 wire \m_blake2.m_hash256.m_matrix[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][6] ;
 wire \m_blake2.m_hash256.m_matrix[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][7] ;
 wire \m_blake2.m_hash256.m_matrix[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][8] ;
 wire \m_blake2.m_hash256.m_matrix[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[8][9] ;
 wire \m_blake2.m_hash256.m_matrix[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][0] ;
 wire \m_blake2.m_hash256.m_matrix[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][10] ;
 wire \m_blake2.m_hash256.m_matrix[9][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][11] ;
 wire \m_blake2.m_hash256.m_matrix[9][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][12] ;
 wire \m_blake2.m_hash256.m_matrix[9][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][13] ;
 wire \m_blake2.m_hash256.m_matrix[9][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][14] ;
 wire \m_blake2.m_hash256.m_matrix[9][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][15] ;
 wire \m_blake2.m_hash256.m_matrix[9][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][16] ;
 wire \m_blake2.m_hash256.m_matrix[9][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][17] ;
 wire \m_blake2.m_hash256.m_matrix[9][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][18] ;
 wire \m_blake2.m_hash256.m_matrix[9][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][19] ;
 wire \m_blake2.m_hash256.m_matrix[9][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][1] ;
 wire \m_blake2.m_hash256.m_matrix[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][20] ;
 wire \m_blake2.m_hash256.m_matrix[9][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][21] ;
 wire \m_blake2.m_hash256.m_matrix[9][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][22] ;
 wire \m_blake2.m_hash256.m_matrix[9][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][23] ;
 wire \m_blake2.m_hash256.m_matrix[9][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][24] ;
 wire \m_blake2.m_hash256.m_matrix[9][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][25] ;
 wire \m_blake2.m_hash256.m_matrix[9][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][26] ;
 wire \m_blake2.m_hash256.m_matrix[9][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][27] ;
 wire \m_blake2.m_hash256.m_matrix[9][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][28] ;
 wire \m_blake2.m_hash256.m_matrix[9][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][29] ;
 wire \m_blake2.m_hash256.m_matrix[9][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][2] ;
 wire \m_blake2.m_hash256.m_matrix[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][30] ;
 wire \m_blake2.m_hash256.m_matrix[9][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][31] ;
 wire \m_blake2.m_hash256.m_matrix[9][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][3] ;
 wire \m_blake2.m_hash256.m_matrix[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][4] ;
 wire \m_blake2.m_hash256.m_matrix[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][5] ;
 wire \m_blake2.m_hash256.m_matrix[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][6] ;
 wire \m_blake2.m_hash256.m_matrix[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][7] ;
 wire \m_blake2.m_hash256.m_matrix[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][8] ;
 wire \m_blake2.m_hash256.m_matrix[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.m_matrix[9][9] ;
 wire \m_blake2.m_hash256.m_matrix[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.res_cnt_q[0] ;
 wire \m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.res_cnt_q[1] ;
 wire \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_blake2.m_hash256.res_cnt_q[2] ;
 wire \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A_X ;
 wire \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.res_cnt_q[3] ;
 wire \m_blake2.m_hash256.res_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.res_cnt_q[4] ;
 wire \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.res_cnt_q[5] ;
 wire \m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.round_q[0] ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_1_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_B1 ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_B_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_A ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_D ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_A ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_C ;
 wire \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1] ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1 ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_1_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1 ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_2_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_3_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o211a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[2] ;
 wire \m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[3] ;
 wire \m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[4] ;
 wire \m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[5] ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_1_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_D ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nand4_2_C_Y ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ;
 wire \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.round_q[6] ;
 wire \m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[7] ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_B ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_A ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_B ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a221o_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_B2_X ;
 wire \m_blake2.m_hash256.round_q[8] ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_A ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_C ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_C ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_C ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o31a_2_A3_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_2_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.round_q[9] ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_A2 ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X_sky130_fd_sc_hd__o21a_2_A2_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X_sky130_fd_sc_hd__o31a_2_A3_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_A2 ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_B1 ;
 wire \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.shift_hash_q ;
 wire \m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1 ;
 wire \m_blake2.m_hash256.slow_output_q ;
 wire \m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][0] ;
 wire \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21oi_2_B1_Y ;
 wire \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.v_q[0][10] ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][11] ;
 wire \m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][12] ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][13] ;
 wire \m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][14] ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][15] ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][16] ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_A2 ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][17] ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][18] ;
 wire \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][19] ;
 wire \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][1] ;
 wire \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][20] ;
 wire \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][21] ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][22] ;
 wire \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][23] ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][24] ;
 wire \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ;
 wire \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][25] ;
 wire \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][26] ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2 ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_X ;
 wire \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][27] ;
 wire \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X ;
 wire \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][28] ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_A2 ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][29] ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_B2 ;
 wire \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][2] ;
 wire \m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][30] ;
 wire \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][31] ;
 wire \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][3] ;
 wire \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][4] ;
 wire \m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][5] ;
 wire \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][6] ;
 wire \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][7] ;
 wire \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][8] ;
 wire \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__and2b_2_B_X ;
 wire \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[0][9] ;
 wire \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[10][0] ;
 wire \m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][10] ;
 wire \m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][11] ;
 wire \m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ;
 wire \m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[10][12] ;
 wire \m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][13] ;
 wire \m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][14] ;
 wire \m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[10][15] ;
 wire \m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][16] ;
 wire \m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][17] ;
 wire \m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][18] ;
 wire \m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][19] ;
 wire \m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[10][1] ;
 wire \m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[10][20] ;
 wire \m_blake2.m_hash256.v_q[10][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][21] ;
 wire \m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[10][22] ;
 wire \m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][23] ;
 wire \m_blake2.m_hash256.v_q[10][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][24] ;
 wire \m_blake2.m_hash256.v_q[10][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][25] ;
 wire \m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][26] ;
 wire \m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][27] ;
 wire \m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[10][28] ;
 wire \m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[10][29] ;
 wire \m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][2] ;
 wire \m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][30] ;
 wire \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ;
 wire \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1_Y ;
 wire \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][31] ;
 wire \m_blake2.m_hash256.v_q[10][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][3] ;
 wire \m_blake2.m_hash256.v_q[10][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][4] ;
 wire \m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[10][5] ;
 wire \m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][6] ;
 wire \m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][7] ;
 wire \m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][8] ;
 wire \m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ;
 wire \m_blake2.m_hash256.v_q[10][9] ;
 wire \m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[11][0] ;
 wire \m_blake2.m_hash256.v_q[11][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][10] ;
 wire \m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][11] ;
 wire \m_blake2.m_hash256.v_q[11][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][12] ;
 wire \m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][13] ;
 wire \m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][14] ;
 wire \m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[11][15] ;
 wire \m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][16] ;
 wire \m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][17] ;
 wire \m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][18] ;
 wire \m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][19] ;
 wire \m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[11][1] ;
 wire \m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ;
 wire \m_blake2.m_hash256.v_q[11][20] ;
 wire \m_blake2.m_hash256.v_q[11][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][21] ;
 wire \m_blake2.m_hash256.v_q[11][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][22] ;
 wire \m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][23] ;
 wire \m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][24] ;
 wire \m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][25] ;
 wire \m_blake2.m_hash256.v_q[11][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][26] ;
 wire \m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][27] ;
 wire \m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][28] ;
 wire \m_blake2.m_hash256.v_q[11][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][29] ;
 wire \m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][2] ;
 wire \m_blake2.m_hash256.v_q[11][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][30] ;
 wire \m_blake2.m_hash256.v_q[11][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][31] ;
 wire \m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][3] ;
 wire \m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][4] ;
 wire \m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][5] ;
 wire \m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][6] ;
 wire \m_blake2.m_hash256.v_q[11][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][7] ;
 wire \m_blake2.m_hash256.v_q[11][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][8] ;
 wire \m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[11][9] ;
 wire \m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][0] ;
 wire \m_blake2.m_hash256.v_q[12][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][10] ;
 wire \m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][11] ;
 wire \m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][12] ;
 wire \m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][13] ;
 wire \m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][14] ;
 wire \m_blake2.m_hash256.v_q[12][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][15] ;
 wire \m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][16] ;
 wire \m_blake2.m_hash256.v_q[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][17] ;
 wire \m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][18] ;
 wire \m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[12][19] ;
 wire \m_blake2.m_hash256.v_q[12][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][1] ;
 wire \m_blake2.m_hash256.v_q[12][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][20] ;
 wire \m_blake2.m_hash256.v_q[12][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][21] ;
 wire \m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][22] ;
 wire \m_blake2.m_hash256.v_q[12][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][23] ;
 wire \m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][24] ;
 wire \m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][25] ;
 wire \m_blake2.m_hash256.v_q[12][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][26] ;
 wire \m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][27] ;
 wire \m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][28] ;
 wire \m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][29] ;
 wire \m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][2] ;
 wire \m_blake2.m_hash256.v_q[12][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][30] ;
 wire \m_blake2.m_hash256.v_q[12][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][31] ;
 wire \m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][3] ;
 wire \m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][4] ;
 wire \m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][5] ;
 wire \m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][6] ;
 wire \m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][7] ;
 wire \m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ;
 wire \m_blake2.m_hash256.v_q[12][8] ;
 wire \m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[12][9] ;
 wire \m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][0] ;
 wire \m_blake2.m_hash256.v_q[13][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][10] ;
 wire \m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][11] ;
 wire \m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[13][12] ;
 wire \m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][13] ;
 wire \m_blake2.m_hash256.v_q[13][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][14] ;
 wire \m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ;
 wire \m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][15] ;
 wire \m_blake2.m_hash256.v_q[13][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][16] ;
 wire \m_blake2.m_hash256.v_q[13][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][17] ;
 wire \m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][18] ;
 wire \m_blake2.m_hash256.v_q[13][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][19] ;
 wire \m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][1] ;
 wire \m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][20] ;
 wire \m_blake2.m_hash256.v_q[13][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][21] ;
 wire \m_blake2.m_hash256.v_q[13][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][22] ;
 wire \m_blake2.m_hash256.v_q[13][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][23] ;
 wire \m_blake2.m_hash256.v_q[13][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][24] ;
 wire \m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ;
 wire \m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][25] ;
 wire \m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[13][26] ;
 wire \m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][27] ;
 wire \m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__nor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[13][28] ;
 wire \m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ;
 wire \m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][29] ;
 wire \m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][2] ;
 wire \m_blake2.m_hash256.v_q[13][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][30] ;
 wire \m_blake2.m_hash256.v_q[13][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][31] ;
 wire \m_blake2.m_hash256.v_q[13][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][3] ;
 wire \m_blake2.m_hash256.v_q[13][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][4] ;
 wire \m_blake2.m_hash256.v_q[13][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][5] ;
 wire \m_blake2.m_hash256.v_q[13][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][6] ;
 wire \m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__a221o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][7] ;
 wire \m_blake2.m_hash256.v_q[13][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][8] ;
 wire \m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[13][9] ;
 wire \m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][0] ;
 wire \m_blake2.m_hash256.v_q[14][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][10] ;
 wire \m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][11] ;
 wire \m_blake2.m_hash256.v_q[14][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][12] ;
 wire \m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][13] ;
 wire \m_blake2.m_hash256.v_q[14][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][14] ;
 wire \m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][15] ;
 wire \m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][16] ;
 wire \m_blake2.m_hash256.v_q[14][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][17] ;
 wire \m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][18] ;
 wire \m_blake2.m_hash256.v_q[14][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][19] ;
 wire \m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][1] ;
 wire \m_blake2.m_hash256.v_q[14][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][20] ;
 wire \m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][21] ;
 wire \m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][22] ;
 wire \m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][23] ;
 wire \m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][24] ;
 wire \m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][25] ;
 wire \m_blake2.m_hash256.v_q[14][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][26] ;
 wire \m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][27] ;
 wire \m_blake2.m_hash256.v_q[14][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][28] ;
 wire \m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][29] ;
 wire \m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][2] ;
 wire \m_blake2.m_hash256.v_q[14][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][30] ;
 wire \m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][31] ;
 wire \m_blake2.m_hash256.v_q[14][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][3] ;
 wire \m_blake2.m_hash256.v_q[14][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][4] ;
 wire \m_blake2.m_hash256.v_q[14][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][5] ;
 wire \m_blake2.m_hash256.v_q[14][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][6] ;
 wire \m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][7] ;
 wire \m_blake2.m_hash256.v_q[14][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][8] ;
 wire \m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[14][9] ;
 wire \m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][0] ;
 wire \m_blake2.m_hash256.v_q[15][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][10] ;
 wire \m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][11] ;
 wire \m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][12] ;
 wire \m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][13] ;
 wire \m_blake2.m_hash256.v_q[15][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][14] ;
 wire \m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][15] ;
 wire \m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][16] ;
 wire \m_blake2.m_hash256.v_q[15][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][17] ;
 wire \m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][18] ;
 wire \m_blake2.m_hash256.v_q[15][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][19] ;
 wire \m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][1] ;
 wire \m_blake2.m_hash256.v_q[15][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][20] ;
 wire \m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][21] ;
 wire \m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][22] ;
 wire \m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][23] ;
 wire \m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][24] ;
 wire \m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][25] ;
 wire \m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][26] ;
 wire \m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][27] ;
 wire \m_blake2.m_hash256.v_q[15][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][28] ;
 wire \m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][29] ;
 wire \m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][2] ;
 wire \m_blake2.m_hash256.v_q[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][30] ;
 wire \m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][31] ;
 wire \m_blake2.m_hash256.v_q[15][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][3] ;
 wire \m_blake2.m_hash256.v_q[15][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][4] ;
 wire \m_blake2.m_hash256.v_q[15][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][5] ;
 wire \m_blake2.m_hash256.v_q[15][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][6] ;
 wire \m_blake2.m_hash256.v_q[15][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][7] ;
 wire \m_blake2.m_hash256.v_q[15][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][8] ;
 wire \m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[15][9] ;
 wire \m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ;
 wire \m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][0] ;
 wire \m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][10] ;
 wire \m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__o22a_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][11] ;
 wire \m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][12] ;
 wire \m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][13] ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][14] ;
 wire \m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][15] ;
 wire \m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][16] ;
 wire \m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][17] ;
 wire \m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][18] ;
 wire \m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][19] ;
 wire \m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][1] ;
 wire \m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][20] ;
 wire \m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][21] ;
 wire \m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][22] ;
 wire \m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][23] ;
 wire \m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][24] ;
 wire \m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][25] ;
 wire \m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][26] ;
 wire \m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][27] ;
 wire \m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][28] ;
 wire \m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][29] ;
 wire \m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][2] ;
 wire \m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][30] ;
 wire \m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][31] ;
 wire \m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][3] ;
 wire \m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][4] ;
 wire \m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][5] ;
 wire \m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][6] ;
 wire \m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][7] ;
 wire \m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][8] ;
 wire \m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[1][9] ;
 wire \m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][0] ;
 wire \m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][10] ;
 wire \m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][11] ;
 wire \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][12] ;
 wire \m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][13] ;
 wire \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][14] ;
 wire \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][15] ;
 wire \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][16] ;
 wire \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][17] ;
 wire \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][18] ;
 wire \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][19] ;
 wire \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][1] ;
 wire \m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][20] ;
 wire \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][21] ;
 wire \m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][22] ;
 wire \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][23] ;
 wire \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][24] ;
 wire \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][25] ;
 wire \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][26] ;
 wire \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][27] ;
 wire \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__a211oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][28] ;
 wire \m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][29] ;
 wire \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__a211oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][2] ;
 wire \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][30] ;
 wire \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][31] ;
 wire \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__a211oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][3] ;
 wire \m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][4] ;
 wire \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__a21oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][5] ;
 wire \m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][6] ;
 wire \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][7] ;
 wire \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[2][8] ;
 wire \m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[2][9] ;
 wire \m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][0] ;
 wire \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][10] ;
 wire \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][11] ;
 wire \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_B1 ;
 wire \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][12] ;
 wire \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][13] ;
 wire \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][14] ;
 wire \m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][15] ;
 wire \m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][16] ;
 wire \m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][17] ;
 wire \m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][18] ;
 wire \m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][19] ;
 wire \m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][1] ;
 wire \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][20] ;
 wire \m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][21] ;
 wire \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__a211oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][22] ;
 wire \m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][23] ;
 wire \m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][24] ;
 wire \m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][25] ;
 wire \m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][26] ;
 wire \m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][27] ;
 wire \m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][28] ;
 wire \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][29] ;
 wire \m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][2] ;
 wire \m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][30] ;
 wire \m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][31] ;
 wire \m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][3] ;
 wire \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][4] ;
 wire \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_B1 ;
 wire \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][5] ;
 wire \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__a211o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][6] ;
 wire \m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][7] ;
 wire \m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[3][8] ;
 wire \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__a211oi_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[3][9] ;
 wire \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__a31o_2_A3_X ;
 wire \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__xor2_2_B_X ;
 wire \m_blake2.m_hash256.v_q[4][0] ;
 wire \m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[4][10] ;
 wire \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][11] ;
 wire \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][12] ;
 wire \m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][13] ;
 wire \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][14] ;
 wire \m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][15] ;
 wire \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][16] ;
 wire \m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][17] ;
 wire \m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][18] ;
 wire \m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][19] ;
 wire \m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][1] ;
 wire \m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[4][20] ;
 wire \m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][21] ;
 wire \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][22] ;
 wire \m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][23] ;
 wire \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][24] ;
 wire \m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][25] ;
 wire \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][26] ;
 wire \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][27] ;
 wire \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][28] ;
 wire \m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][29] ;
 wire \m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][2] ;
 wire \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[4][30] ;
 wire \m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][31] ;
 wire \m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][3] ;
 wire \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[4][4] ;
 wire \m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[4][5] ;
 wire \m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[4][6] ;
 wire \m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[4][7] ;
 wire \m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][8] ;
 wire \m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[4][9] ;
 wire \m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][0] ;
 wire \m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][10] ;
 wire \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][11] ;
 wire \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][12] ;
 wire \m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][13] ;
 wire \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][14] ;
 wire \m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][15] ;
 wire \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][16] ;
 wire \m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][17] ;
 wire \m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][18] ;
 wire \m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][19] ;
 wire \m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][1] ;
 wire \m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][20] ;
 wire \m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][21] ;
 wire \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][22] ;
 wire \m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][23] ;
 wire \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][24] ;
 wire \m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][25] ;
 wire \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][26] ;
 wire \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][27] ;
 wire \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][28] ;
 wire \m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][29] ;
 wire \m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][2] ;
 wire \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[5][30] ;
 wire \m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][31] ;
 wire \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__mux2_1_A0_1_X ;
 wire \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][3] ;
 wire \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[5][4] ;
 wire \m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][5] ;
 wire \m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][6] ;
 wire \m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[5][7] ;
 wire \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[5][8] ;
 wire \m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[5][9] ;
 wire \m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][0] ;
 wire \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[6][10] ;
 wire \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][11] ;
 wire \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][12] ;
 wire \m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][13] ;
 wire \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][14] ;
 wire \m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][15] ;
 wire \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][16] ;
 wire \m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][17] ;
 wire \m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][18] ;
 wire \m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][19] ;
 wire \m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][1] ;
 wire \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[6][20] ;
 wire \m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][21] ;
 wire \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][22] ;
 wire \m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][23] ;
 wire \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][24] ;
 wire \m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][25] ;
 wire \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][26] ;
 wire \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][27] ;
 wire \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ;
 wire \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][28] ;
 wire \m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][29] ;
 wire \m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][2] ;
 wire \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][30] ;
 wire \m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][31] ;
 wire \m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][3] ;
 wire \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[6][4] ;
 wire \m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][5] ;
 wire \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[6][6] ;
 wire \m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][7] ;
 wire \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[6][8] ;
 wire \m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[6][9] ;
 wire \m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][0] ;
 wire \m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[7][10] ;
 wire \m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][11] ;
 wire \m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][12] ;
 wire \m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][13] ;
 wire \m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][14] ;
 wire \m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][15] ;
 wire \m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][16] ;
 wire \m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][17] ;
 wire \m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][18] ;
 wire \m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][19] ;
 wire \m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][1] ;
 wire \m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][20] ;
 wire \m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][21] ;
 wire \m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][22] ;
 wire \m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][23] ;
 wire \m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][24] ;
 wire \m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][25] ;
 wire \m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][26] ;
 wire \m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][27] ;
 wire \m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][28] ;
 wire \m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][29] ;
 wire \m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][2] ;
 wire \m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][30] ;
 wire \m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][31] ;
 wire \m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][3] ;
 wire \m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[7][4] ;
 wire \m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[7][5] ;
 wire \m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][6] ;
 wire \m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][7] ;
 wire \m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[7][8] ;
 wire \m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[7][9] ;
 wire \m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[8][0] ;
 wire \m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][10] ;
 wire \m_blake2.m_hash256.v_q[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][11] ;
 wire \m_blake2.m_hash256.v_q[8][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][12] ;
 wire \m_blake2.m_hash256.v_q[8][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][13] ;
 wire \m_blake2.m_hash256.v_q[8][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][14] ;
 wire \m_blake2.m_hash256.v_q[8][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][15] ;
 wire \m_blake2.m_hash256.v_q[8][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][16] ;
 wire \m_blake2.m_hash256.v_q[8][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][17] ;
 wire \m_blake2.m_hash256.v_q[8][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][18] ;
 wire \m_blake2.m_hash256.v_q[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][19] ;
 wire \m_blake2.m_hash256.v_q[8][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][1] ;
 wire \m_blake2.m_hash256.v_q[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][20] ;
 wire \m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][21] ;
 wire \m_blake2.m_hash256.v_q[8][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][22] ;
 wire \m_blake2.m_hash256.v_q[8][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][23] ;
 wire \m_blake2.m_hash256.v_q[8][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][24] ;
 wire \m_blake2.m_hash256.v_q[8][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][25] ;
 wire \m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_blake2.m_hash256.v_q[8][26] ;
 wire \m_blake2.m_hash256.v_q[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][27] ;
 wire \m_blake2.m_hash256.v_q[8][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][28] ;
 wire \m_blake2.m_hash256.v_q[8][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][29] ;
 wire \m_blake2.m_hash256.v_q[8][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][2] ;
 wire \m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][30] ;
 wire \m_blake2.m_hash256.v_q[8][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][31] ;
 wire \m_blake2.m_hash256.v_q[8][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][3] ;
 wire \m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ;
 wire \m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][4] ;
 wire \m_blake2.m_hash256.v_q[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][5] ;
 wire \m_blake2.m_hash256.v_q[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][6] ;
 wire \m_blake2.m_hash256.v_q[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][7] ;
 wire \m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][8] ;
 wire \m_blake2.m_hash256.v_q[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[8][9] ;
 wire \m_blake2.m_hash256.v_q[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][0] ;
 wire \m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][10] ;
 wire \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][11] ;
 wire \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][12] ;
 wire \m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][13] ;
 wire \m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][14] ;
 wire \m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][15] ;
 wire \m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][16] ;
 wire \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__o21a_2_A1_X ;
 wire \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][17] ;
 wire \m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][18] ;
 wire \m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][19] ;
 wire \m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][1] ;
 wire \m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][20] ;
 wire \m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][21] ;
 wire \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][22] ;
 wire \m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][23] ;
 wire \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__a22o_2_B1_X ;
 wire \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][24] ;
 wire \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][25] ;
 wire \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A ;
 wire \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_X ;
 wire \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][26] ;
 wire \m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][27] ;
 wire \m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][28] ;
 wire \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][29] ;
 wire \m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][2] ;
 wire \m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][30] ;
 wire \m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][31] ;
 wire \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][3] ;
 wire \m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][4] ;
 wire \m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][5] ;
 wire \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ;
 wire \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_Y ;
 wire \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ;
 wire \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_A ;
 wire \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][6] ;
 wire \m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][7] ;
 wire \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][8] ;
 wire \m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_blake2.m_hash256.v_q[9][9] ;
 wire \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_io.cmd[1] ;
 wire \m_io.cmd[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.cmd[2] ;
 wire \m_io.cmd[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.cmd[2]_sky130_fd_sc_hd__o21ai_2_A1_Y ;
 wire \m_io.cmd[4] ;
 wire \m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_io.cmd[5] ;
 wire \m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B ;
 wire \m_io.data_v_early ;
 wire \m_io.data_v_early_sky130_fd_sc_hd__a21oi_2_A2_Y ;
 wire \m_io.data_v_early_sky130_fd_sc_hd__and3_2_C_X ;
 wire \m_io.en_q ;
 wire \m_io.en_q_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.hash_v_o ;
 wire \m_io.m_block_data.data_cnt_q[0] ;
 wire \m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_io.m_block_data.data_cnt_q[1] ;
 wire \m_io.m_block_data.data_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_block_data.data_cnt_q[2] ;
 wire \m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_io.m_block_data.data_cnt_q[3] ;
 wire \m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_B ;
 wire \m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_C ;
 wire \m_io.m_block_data.data_cnt_q[4] ;
 wire \m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B ;
 wire \m_io.m_block_data.data_cnt_q[5] ;
 wire \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_D ;
 wire \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_X ;
 wire \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_B ;
 wire \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_io.m_config.cfg_cnt_q[0] ;
 wire \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A ;
 wire \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ;
 wire \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_B ;
 wire \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C ;
 wire \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B ;
 wire \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_io.m_config.cfg_cnt_q[1] ;
 wire \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N ;
 wire \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ;
 wire \m_io.m_config.cfg_cnt_q[2] ;
 wire \m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_io.m_config.cfg_cnt_q[3] ;
 wire \m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire \m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__nand3_2_C_Y ;
 wire \m_io.m_config.data_i[0] ;
 wire \m_io.m_config.data_i[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.data_i[1] ;
 wire \m_io.m_config.data_i[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.data_i[2] ;
 wire \m_io.m_config.data_i[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.data_i[3] ;
 wire \m_io.m_config.data_i[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.data_i[4] ;
 wire \m_io.m_config.data_i[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.data_i[5] ;
 wire \m_io.m_config.data_i[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.data_i[6] ;
 wire \m_io.m_config.data_i[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.data_i[7] ;
 wire \m_io.m_config.data_i[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.kk_q[0] ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__mux2_1_A1_X ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ;
 wire \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ;
 wire \m_io.m_config.kk_q[1] ;
 wire \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_io.m_config.kk_q[2] ;
 wire \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_io.m_config.kk_q[3] ;
 wire \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X ;
 wire \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ;
 wire \m_io.m_config.kk_q[4] ;
 wire \m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1_X ;
 wire \m_io.m_config.kk_q[5] ;
 wire \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ;
 wire \m_io.m_config.ll_q[0] ;
 wire \m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[10] ;
 wire \m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[11] ;
 wire \m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[12] ;
 wire \m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[13] ;
 wire \m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[14] ;
 wire \m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[15] ;
 wire \m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[16] ;
 wire \m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[17] ;
 wire \m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[18] ;
 wire \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ;
 wire \m_io.m_config.ll_q[19] ;
 wire \m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[1] ;
 wire \m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[20] ;
 wire \m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[21] ;
 wire \m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[22] ;
 wire \m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[23] ;
 wire \m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[24] ;
 wire \m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[25] ;
 wire \m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[26] ;
 wire \m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[27] ;
 wire \m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[28] ;
 wire \m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[29] ;
 wire \m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[2] ;
 wire \m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[30] ;
 wire \m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[31] ;
 wire \m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[32] ;
 wire \m_io.m_config.ll_q[32]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[33] ;
 wire \m_io.m_config.ll_q[33]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[34] ;
 wire \m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[35] ;
 wire \m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[36] ;
 wire \m_io.m_config.ll_q[36]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[37] ;
 wire \m_io.m_config.ll_q[37]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[38] ;
 wire \m_io.m_config.ll_q[38]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[39] ;
 wire \m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[3] ;
 wire \m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[40] ;
 wire \m_io.m_config.ll_q[40]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[41] ;
 wire \m_io.m_config.ll_q[41]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[42] ;
 wire \m_io.m_config.ll_q[42]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[43] ;
 wire \m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[44] ;
 wire \m_io.m_config.ll_q[44]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[45] ;
 wire \m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[46] ;
 wire \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ;
 wire \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ;
 wire \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ;
 wire \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ;
 wire \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[47] ;
 wire \m_io.m_config.ll_q[47]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[48] ;
 wire \m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[49] ;
 wire \m_io.m_config.ll_q[49]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[4] ;
 wire \m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[50] ;
 wire \m_io.m_config.ll_q[50]_sky130_fd_sc_hd__a22o_2_B2_X ;
 wire \m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[51] ;
 wire \m_io.m_config.ll_q[51]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[52] ;
 wire \m_io.m_config.ll_q[52]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[53] ;
 wire \m_io.m_config.ll_q[53]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[54] ;
 wire \m_io.m_config.ll_q[54]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[55] ;
 wire \m_io.m_config.ll_q[55]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[56] ;
 wire \m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[57] ;
 wire \m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[58] ;
 wire \m_io.m_config.ll_q[58]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[59] ;
 wire \m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[5] ;
 wire \m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[60] ;
 wire \m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[61] ;
 wire \m_io.m_config.ll_q[61]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[62] ;
 wire \m_io.m_config.ll_q[62]_sky130_fd_sc_hd__and3_2_A_X ;
 wire \m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[63] ;
 wire \m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[6] ;
 wire \m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[7] ;
 wire \m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[8] ;
 wire \m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.ll_q[9] ;
 wire \m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.nn_q[0] ;
 wire \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ;
 wire \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__or2_2_A_B ;
 wire \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A_X ;
 wire \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X ;
 wire \m_io.m_config.nn_q[1] ;
 wire \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_io.m_config.nn_q[2] ;
 wire \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_io.m_config.nn_q[3] ;
 wire \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ;
 wire \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ;
 wire \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ;
 wire \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_io.m_config.nn_q[4] ;
 wire \m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.nn_q[5] ;
 wire \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ;
 wire \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y ;
 wire \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y ;
 wire \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A_B ;
 wire \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A_C ;
 wire \m_io.m_config.valid_i ;
 wire \m_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q_D ;
 wire \m_io.ready_v_o ;
 wire \m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1 ;
 wire net628;
 wire net627;
 wire net626;
 wire clknet_leaf_0_clk;
 wire net625;
 wire net624;
 wire net623;
 wire net635;
 wire net634;
 wire net633;
 wire net632;
 wire net631;
 wire net630;
 wire net629;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_A2;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_B1;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X_B1;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X_B1;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2;
 wire uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_0_clk;
 wire clknet_3_0_0_clk;
 wire clknet_3_1_0_clk;
 wire clknet_3_2_0_clk;
 wire clknet_3_3_0_clk;
 wire clknet_3_4_0_clk;
 wire clknet_3_5_0_clk;
 wire clknet_3_6_0_clk;
 wire clknet_3_7_0_clk;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;

 sky130_fd_sc_hd__a22o_1 block_first_sky130_fd_sc_hd__a22o_2_B2 (.A1(net485),
    .A2(block_last_sky130_fd_sc_hd__a22o_2_B2_A2),
    .B1(block_last_sky130_fd_sc_hd__a22o_2_B2_B1),
    .B2(net648),
    .X(\m_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a32o_1 block_first_sky130_fd_sc_hd__a32o_2_B2 (.A1(block_first_sky130_fd_sc_hd__a32o_2_B2_A1),
    .A2(\m_io.cmd[1] ),
    .A3(\m_io.m_config.valid_i ),
    .B1(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_X ),
    .B2(block_first),
    .X(block_first_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B));
 sky130_fd_sc_hd__clkinv_2 block_first_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__inv_2_Y (.A(\m_io.cmd[2] ),
    .Y(block_first_sky130_fd_sc_hd__a32o_2_B2_A1));
 sky130_fd_sc_hd__dfxtp_1 block_first_sky130_fd_sc_hd__dfxtp_2_Q (.CLK(clknet_leaf_21_clk),
    .D(block_first_sky130_fd_sc_hd__dfxtp_2_Q_D),
    .Q(block_first));
 sky130_fd_sc_hd__and2_1 block_first_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X (.A(net610),
    .B(block_first_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B),
    .X(block_first_sky130_fd_sc_hd__dfxtp_2_Q_D));
 sky130_fd_sc_hd__a22o_1 block_last_sky130_fd_sc_hd__a22o_2_B2 (.A1(net463),
    .A2(block_last_sky130_fd_sc_hd__a22o_2_B2_A2),
    .B1(block_last_sky130_fd_sc_hd__a22o_2_B2_B1),
    .B2(net655),
    .X(\m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 block_last_sky130_fd_sc_hd__a22o_2_B2_B1_sky130_fd_sc_hd__nor2_2_Y (.A(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(block_last_sky130_fd_sc_hd__a22o_2_B2_A2),
    .Y(block_last_sky130_fd_sc_hd__a22o_2_B2_B1));
 sky130_fd_sc_hd__a32o_1 block_last_sky130_fd_sc_hd__a32o_2_B2 (.A1(\m_io.cmd[2] ),
    .A2(\m_io.cmd[1] ),
    .A3(\m_io.m_config.valid_i ),
    .B1(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_X ),
    .B2(block_last),
    .X(block_last_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B));
 sky130_fd_sc_hd__dfxtp_1 block_last_sky130_fd_sc_hd__dfxtp_2_Q (.CLK(clknet_leaf_21_clk),
    .D(block_last_sky130_fd_sc_hd__dfxtp_2_Q_D),
    .Q(block_last));
 sky130_fd_sc_hd__and2_1 block_last_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X (.A(net610),
    .B(block_last_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B),
    .X(block_last_sky130_fd_sc_hd__dfxtp_2_Q_D));
 sky130_fd_sc_hd__dfxtp_1 \data[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\data[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[0] ));
 sky130_fd_sc_hd__mux2_1 \data[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[0] ),
    .A1(net644),
    .S(net308),
    .X(\data[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[0]_sky130_fd_sc_hd__mux2_1_A1  (.A0(net646),
    .A1(net644),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[15][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \data[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\data[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[1] ));
 sky130_fd_sc_hd__mux2_1 \data[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[1] ),
    .A1(net647),
    .S(net308),
    .X(\data[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[1]_sky130_fd_sc_hd__mux2_1_A1  (.A0(net649),
    .A1(net647),
    .S(net589),
    .X(\m_blake2.m_hash256.m_matrix[15][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \data[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\data[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[2] ));
 sky130_fd_sc_hd__mux2_1 \data[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[2] ),
    .A1(net650),
    .S(net308),
    .X(\data[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[2]_sky130_fd_sc_hd__mux2_1_A1  (.A0(net651),
    .A1(net650),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[15][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \data[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\data[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[3] ));
 sky130_fd_sc_hd__mux2_1 \data[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[3] ),
    .A1(net642),
    .S(net308),
    .X(\data[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[3]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_matrix[15][27] ),
    .A1(net642),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[15][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \data[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\data[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[4] ));
 sky130_fd_sc_hd__mux2_1 \data[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[4] ),
    .A1(net814),
    .S(net308),
    .X(\data[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[4]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_matrix[15][28] ),
    .A1(net814),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[15][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \data[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\data[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[5] ));
 sky130_fd_sc_hd__mux2_1 \data[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[5] ),
    .A1(net1682),
    .S(net308),
    .X(\data[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[5]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_matrix[15][29] ),
    .A1(net1682),
    .S(net550),
    .X(\m_blake2.m_hash256.m_matrix[15][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \data[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\data[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[6] ));
 sky130_fd_sc_hd__mux2_1 \data[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[6] ),
    .A1(net834),
    .S(\m_io.cmd[2]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .X(\data[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[6]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_matrix[15][30] ),
    .A1(net834),
    .S(net579),
    .X(\m_blake2.m_hash256.m_matrix[15][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \data[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\data[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\data[7] ));
 sky130_fd_sc_hd__mux2_1 \data[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.m_config.data_i[7] ),
    .A1(net874),
    .S(net308),
    .X(\data[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \data[7]_sky130_fd_sc_hd__mux2_1_A1  (.A0(net935),
    .A1(net874),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[15][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and4_1 \data_idx[0]_sky130_fd_sc_hd__and4_2_B  (.A(net599),
    .B(\data_idx[0] ),
    .C(\data_idx[1] ),
    .D(\data_idx[2] ),
    .X(\data_idx[0]_sky130_fd_sc_hd__and4_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \data_idx[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(net640),
    .Q(\data_idx[0] ));
 sky130_fd_sc_hd__dfxtp_1 \data_idx[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(net636),
    .Q(\data_idx[1] ));
 sky130_fd_sc_hd__dfxtp_1 \data_idx[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(net641),
    .Q(\data_idx[2] ));
 sky130_fd_sc_hd__and4_1 \data_idx[3]_sky130_fd_sc_hd__and4_2_A  (.A(\data_idx[3] ),
    .B(\data_idx[4] ),
    .C(\data_idx[5] ),
    .D(\data_idx[0]_sky130_fd_sc_hd__and4_2_B_X ),
    .X(\data_idx[3]_sky130_fd_sc_hd__and4_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \data_idx[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(net637),
    .Q(\data_idx[3] ));
 sky130_fd_sc_hd__dfxtp_1 \data_idx[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(net639),
    .Q(\data_idx[4] ));
 sky130_fd_sc_hd__dfxtp_1 \data_idx[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(net638),
    .Q(\data_idx[5] ));
 sky130_fd_sc_hd__dfxtp_1 data_v_sky130_fd_sc_hd__dfxtp_2_Q (.CLK(clknet_leaf_20_clk),
    .D(\m_io.data_v_early ),
    .Q(data_v));
 sky130_fd_sc_hd__or2_1 ena_sky130_fd_sc_hd__or2_2_B (.A(ena_sky130_fd_sc_hd__or2_2_B_A),
    .B(net1),
    .X(\m_io.en_q_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 ena_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__inv_2_Y (.A(net609),
    .Y(ena_sky130_fd_sc_hd__or2_2_B_A));
 sky130_fd_sc_hd__dfxtp_2 \hash[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[0] ));
 sky130_fd_sc_hd__mux2_1 \hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[0] ),
    .S(net309),
    .X(\hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \hash[0]_sky130_fd_sc_hd__or2_2_B  (.A(net483),
    .B(\hash[0] ),
    .X(\hash[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and3_1 \hash[0]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C  (.A(net402),
    .B(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\hash[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\hash[0]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \hash[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\hash[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[1] ));
 sky130_fd_sc_hd__mux2_1 \hash[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[1] ),
    .S(net316),
    .X(\hash[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_2 \hash[1]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A1(\hash[1] ),
    .S(net430),
    .X(\hash[1]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \hash[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\hash[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[2] ));
 sky130_fd_sc_hd__mux2_1 \hash[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[2] ),
    .S(net316),
    .X(\hash[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \hash[2]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A1(\hash[2] ),
    .S(net430),
    .X(\hash[2]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__a221oi_1 \hash[2]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2  (.A1(net401),
    .A2(\hash[2]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .B1(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net285),
    .C1(net345),
    .Y(\hash[2]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_2 \hash[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[3] ));
 sky130_fd_sc_hd__mux2_1 \hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[3] ),
    .S(net320),
    .X(\hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_4 \hash[3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\hash[3] ),
    .A1(\m_io.m_config.nn_q[3] ),
    .S(net485),
    .X(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__dfxtp_2 \hash[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[4] ));
 sky130_fd_sc_hd__mux2_1 \hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[4] ),
    .S(net309),
    .X(\hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_4 \hash[4]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\hash[4] ),
    .A1(\m_io.m_config.nn_q[4] ),
    .S(net485),
    .X(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nand2_1 \hash[4]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B  (.A(net403),
    .B(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .Y(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and3_1 \hash[4]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .C(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_B1 ));
 sky130_fd_sc_hd__dfxtp_2 \hash[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[5] ));
 sky130_fd_sc_hd__mux2_1 \hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[5] ),
    .S(net314),
    .X(\hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_4 \hash[5]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A1(\hash[5] ),
    .S(net428),
    .X(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__dfxtp_4 \hash[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[6] ));
 sky130_fd_sc_hd__mux2_1 \hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[6] ),
    .S(net335),
    .X(\hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \hash[6]_sky130_fd_sc_hd__or2_2_B  (.A(net500),
    .B(\hash[6] ),
    .X(\hash[6]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \hash[7]_sky130_fd_sc_hd__and2_2_B  (.A(net442),
    .B(\hash[7] ),
    .X(\hash[7]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_4 \hash[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\hash[7] ));
 sky130_fd_sc_hd__mux2_1 \hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\hash[7] ),
    .S(net335),
    .X(\hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a211o_1 hash_v_sky130_fd_sc_hd__a211o_2_X (.A1(net463),
    .A2(\m_blake2.m_hash256.fsm_q[5] ),
    .B1(net656),
    .C1(net478),
    .X(hash_v));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[0] ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_A2 ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2 ),
    .B1(net427),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[0] ),
    .B(\m_blake2.m_hash256.f_finished ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2 ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[8] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[9] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[10] ),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[10] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(net1880),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[8] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[9] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[11] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[11] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[11] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(net422),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[12] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(net426),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[11] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[12] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[11] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[12] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[13] ),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[13] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(net1016),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net426),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[11] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[12] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[14] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[14] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[14] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[15] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(net425),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[14] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[15] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[14] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[15] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[16] ),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[16] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(net1149),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net425),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[14] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[15] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[17] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[17] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[17] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(net422),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[18] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(net426),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[17] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[18] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[17] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[18] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[19] ),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[19] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[19] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net426),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[17] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[18] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[0] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[1] ),
    .C(net445),
    .D(\m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[1] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[1] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_A2 ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_X ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[20] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[20] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[20] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[21] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(net426),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[20] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[21] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[20] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[21] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[22] ),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[22] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__and4_2_C_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(net1687),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[20] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[21] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[23] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[23] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(net425),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[23] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[24] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[24] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(net1151),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net425),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[23] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[22]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[25] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[25] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[25] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[26] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[26] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[26] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[26] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[25] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[24]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[27] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[26] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[27] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[27] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net423),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[28] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[28] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[28] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[29] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[29] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[29] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[2] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[2] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[2] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_X ),
    .B1(net427),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[28] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[29] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[30] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[29] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[30] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[30] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net423),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[31] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[31] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[31] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net425),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[32] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[32] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[32] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[31] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[32] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[33] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[32] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[33] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[33] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net425),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[34] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[34] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net1895),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net426),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[35] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[35] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[35] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net422),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[34] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[35] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[36] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[35] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[36] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[36] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net426),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[37] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[37] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[37] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net425),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[38] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[38] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[38] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[37] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[38] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[39] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[38] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[39] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[39] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net425),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[3] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net1859),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1(net427),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[40] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[40] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net1643),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net424),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[41] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[41] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[41] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[40] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[41] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[42] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[41] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[42] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[42] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net424),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[43] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[43] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[43] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net426),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[44] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(net1796),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[44] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[43] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[44] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[45] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[44] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[45] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[45] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net426),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[46] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[46] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net1795),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net425),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[47] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[47] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[47] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net422),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[46] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[47] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[48] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[47] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[48] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[48] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net425),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[49] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[49] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[49] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net424),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[2] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[3] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[4] ),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[4] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(net1464),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net427),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[2] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[3] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[50] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(net1889),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[50] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[49] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[50] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[51] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[50] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[51] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[51] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net424),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[52] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[52] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_C ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[52] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net424),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[53] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[53] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[53] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[52] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[53] ),
    .A3(\m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[54] ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[53] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[54] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[54] ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(net424),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[55] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net1890),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net426),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[55] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[56] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[56] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(net1465),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net427),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[55] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[54]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[57] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(net421),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(net795),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[57] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__o21a_2_A1  (.A1(net794),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__and3_2_B_X ),
    .B1(\m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[5] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[5] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[5] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(net424),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[6] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net1896),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[5] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[6] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[7] ),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[7] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_X ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[7] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[5] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[6] ),
    .C(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[8] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[8] ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_X ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[8] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_X ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.block_idx_plus_one_q[9] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[10]_sky130_fd_sc_hd__o21ai_2_A1_A2 ),
    .B(\m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[9] ),
    .A2(\m_blake2.m_hash256.block_idx_plus_one_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1(net423),
    .Y(\m_blake2.m_hash256.block_idx_plus_one_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.f_finished_q_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.f_finished ),
    .Q(\m_blake2.m_hash256.f_finished_q ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X  (.A(net445),
    .B(\m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.f_finished ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_A_sky130_fd_sc_hd__and3_2_X  (.A(net467),
    .B(net469),
    .C(net474),
    .X(\m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_A ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.block_idx_plus_one_q[0] ),
    .B(net445),
    .C(\m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_A2 ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and4_2_X  (.A(net449),
    .B(\m_blake2.m_hash256.g_idx_next[2] ),
    .C(\m_blake2.m_hash256.g_idx_next[1] ),
    .D(\m_blake2.m_hash256.g_idx_next[0] ),
    .X(\m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.first_block_q ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__inv_2_A  (.A(net495),
    .Y(\hash[7]_sky130_fd_sc_hd__and2_2_B_A ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.fsm_q[0] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.fsm_q[0] ),
    .A2(\m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .B1(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net478),
    .C1(ena_sky130_fd_sc_hd__or2_2_B_A),
    .X(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__nor2_2_B  (.A(net478),
    .B(\m_blake2.m_hash256.fsm_q[0] ),
    .Y(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__or2_4 \m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B  (.A(net478),
    .B(\m_blake2.m_hash256.fsm_q[0] ),
    .X(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.fsm_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.fsm_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.fsm_q[1] ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.fsm_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and4_2_X  (.A(net610),
    .B(net463),
    .C(net1903),
    .D(\m_blake2.m_hash256.fsm_q[5] ),
    .X(\m_blake2.m_hash256.fsm_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.fsm_q[2] ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X  (.A1(net610),
    .A2(\m_blake2.m_hash256.fsm_q[3] ),
    .A3(\data_idx[3]_sky130_fd_sc_hd__and4_2_A_X ),
    .B1(\m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X_B1 ),
    .X(\m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.f_finished ),
    .B(net482),
    .C(net611),
    .X(\m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.fsm_q[3] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\data_idx[3]_sky130_fd_sc_hd__and4_2_A_X ),
    .A2_N(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(net611),
    .B2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2 ),
    .X(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__nand2_2_Y  (.A(net610),
    .B(\m_blake2.m_hash256.fsm_q[3] ),
    .Y(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.fsm_q[5] ),
    .B1(\m_blake2.m_hash256.fsm_q[0] ),
    .B2(net606),
    .X(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2 ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__inv_2_Y  (.A(net463),
    .Y(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1 ));
 sky130_fd_sc_hd__nand2_8 \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1 ),
    .B(net368),
    .Y(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1 ),
    .B(net343),
    .Y(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.fsm_q[4] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(net656),
    .A2(\m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2 ),
    .B1(net611),
    .X(\m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a32o_2_X  (.A1(net463),
    .A2(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A_Y ),
    .A3(\m_blake2.m_hash256.fsm_q[5] ),
    .B1(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__inv_2_Y_A ),
    .B2(net478),
    .X(\m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.fsm_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.fsm_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.fsm_q[5] ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.fsm_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net610),
    .B(net482),
    .C(\m_blake2.m_hash256.f_finished ),
    .X(\m_blake2.m_hash256.fsm_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor3b_1 \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__nor3b_2_C_N  (.A(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2 ),
    .C_N(\m_blake2.m_hash256.g_b[0] ),
    .Y(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[0] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net347),
    .A2_N(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net256),
    .X(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X  (.A1_N(net188),
    .A2_N(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(net274),
    .B2(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net347),
    .A2(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net177),
    .X(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net347),
    .B(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.v_q[4][0] ),
    .A2(net347),
    .B1(net181),
    .X(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[10] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net181),
    .A2(\m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .B(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .B(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .X(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[11] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net184),
    .A2(\m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net102),
    .B2(\m_blake2.m_hash256.m_matrix[0][11] ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][11] ),
    .A2(net127),
    .B1(net114),
    .B2(\m_blake2.m_hash256.m_matrix[5][11] ),
    .C1(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][11] ),
    .A2(net131),
    .B1(net147),
    .B2(\m_blake2.m_hash256.m_matrix[10][11] ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][11] ),
    .A2(net136),
    .B1(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][11] ),
    .A2(net135),
    .B1(net118),
    .B2(\m_blake2.m_hash256.m_matrix[13][11] ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][11] ),
    .A2(net87),
    .B1(net90),
    .B2(\m_blake2.m_hash256.m_matrix[14][11] ),
    .C1(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][11] ),
    .A2(net108),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][11] ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][11] ),
    .A2(net140),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][11] ),
    .C1(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][11] ),
    .A2(net99),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][11] ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[12] ),
    .B(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2  (.A1(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .A2(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__o22a_4 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net182),
    .X(\m_blake2.m_hash256.g_b[12] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net258),
    .A2(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net394),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net199),
    .A2(\m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net191),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net358),
    .A2(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net179),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][12] ),
    .A1(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net395),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[12] ),
    .B(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[13] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__o21ai_4 \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net182),
    .A2(\m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[14] ),
    .B(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A2  (.A1(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ),
    .A2(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ),
    .B(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net183),
    .X(\m_blake2.m_hash256.g_b[14] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net258),
    .A2(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net382),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .A2(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net353),
    .A2(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net180),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][14] ),
    .A1(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net382),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[14] ),
    .B(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[15] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__nor3_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B ));
 sky130_fd_sc_hd__o21ai_4 \m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net182),
    .A2(\m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[16] ),
    .B(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2  (.A1(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1_N(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B  (.A(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X ),
    .C_N(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_b[16] ),
    .B(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__nor3_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net181),
    .X(\m_blake2.m_hash256.g_b[16] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X  (.A(net349),
    .B(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(net256),
    .A2(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net376),
    .C1(net178),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net196),
    .A2(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net188),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][16] ),
    .A1(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net376),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[17] ),
    .B(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net181),
    .X(\m_blake2.m_hash256.g_b[17] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net255),
    .A2(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net367),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net195),
    .A2(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net187),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net345),
    .A2(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net177),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][17] ),
    .A1(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net371),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[17] ),
    .B(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.g_b[18] ),
    .A2(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1 ),
    .Y(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B ),
    .C(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][18] ),
    .B(net102),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_A ));
 sky130_fd_sc_hd__or4_2 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X  (.A(net107),
    .B(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][18] ),
    .A2(net123),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][18] ),
    .C1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][18] ),
    .A2(net127),
    .B1(net147),
    .B2(\m_blake2.m_hash256.m_matrix[10][18] ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][18] ),
    .A2(net91),
    .B1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][18] ),
    .A2(net131),
    .B1(net139),
    .B2(\m_blake2.m_hash256.m_matrix[2][18] ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][18] ),
    .A2(net111),
    .B1(net115),
    .B2(\m_blake2.m_hash256.m_matrix[5][18] ),
    .C1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][18] ),
    .A2(net142),
    .B1(net95),
    .B2(\m_blake2.m_hash256.m_matrix[12][18] ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][18] ),
    .A2(net87),
    .B1(net119),
    .B2(\m_blake2.m_hash256.m_matrix[13][18] ),
    .C1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][18] ),
    .A2(net135),
    .B1(net99),
    .B2(\m_blake2.m_hash256.m_matrix[6][18] ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net181),
    .X(\m_blake2.m_hash256.g_b[18] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net256),
    .A2(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net373),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net196),
    .A2(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net188),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net347),
    .A2(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net177),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][18] ),
    .A1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net374),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[18] ),
    .B(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1 ),
    .B(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .A2(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1 ),
    .A2(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2 ),
    .B1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B2(\m_blake2.m_hash256.g_b[19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_X ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][19] ),
    .A2(net101),
    .B1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][19] ),
    .A2(net86),
    .B1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net107),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][19] ),
    .A2(net126),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][19] ),
    .A2(net111),
    .B1(net131),
    .B2(\m_blake2.m_hash256.m_matrix[8][19] ),
    .C1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][19] ),
    .A2(net91),
    .B1(net135),
    .B2(\m_blake2.m_hash256.m_matrix[3][19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][19] ),
    .A2(net116),
    .B1(net99),
    .B2(\m_blake2.m_hash256.m_matrix[6][19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][19] ),
    .A2(net136),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][19] ),
    .A2(net115),
    .B1(net141),
    .B2(\m_blake2.m_hash256.m_matrix[1][19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][19] ),
    .A2(net121),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21bo_2_X_B1_N ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net181),
    .X(\m_blake2.m_hash256.g_b[19] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net255),
    .A2(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net373),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net196),
    .A2(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net188),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net348),
    .A2(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net178),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][19] ),
    .A1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net375),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[19] ),
    .B(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1 ),
    .B(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2 ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a221o_2_C1  (.A1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .A2(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__inv_2_A_Y ),
    .C1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a221o_2_C1_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[1] ),
    .B(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[1] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net345),
    .A2_N(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net255),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X  (.A1_N(net187),
    .A2_N(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net274),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net345),
    .A2(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net177),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net345),
    .B(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.v_q[4][1] ),
    .A2(net345),
    .B1(net181),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[1] ),
    .B(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__or3b_2_X_C_N ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[20] ),
    .B(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__o32ai_4 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y  (.A1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1 ),
    .A2(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2 ),
    .A3(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3 ),
    .B1(net100),
    .B2(\m_blake2.m_hash256.m_matrix[0][20] ),
    .Y(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][20] ),
    .A2(net144),
    .B1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net104),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][20] ),
    .A2(net128),
    .B1(net96),
    .B2(\m_blake2.m_hash256.m_matrix[6][20] ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][20] ),
    .A2(net108),
    .B1(net136),
    .B2(\m_blake2.m_hash256.m_matrix[2][20] ),
    .C1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][20] ),
    .A2(net92),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][20] ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][20] ),
    .A2(net132),
    .B1(net140),
    .B2(\m_blake2.m_hash256.m_matrix[1][20] ),
    .C1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][20] ),
    .A2(net84),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][20] ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][20] ),
    .A2(net112),
    .B1(net116),
    .B2(\m_blake2.m_hash256.m_matrix[13][20] ),
    .C1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][20] ),
    .A2(net124),
    .B1(net88),
    .B2(\m_blake2.m_hash256.m_matrix[14][20] ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B  (.A(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ),
    .B(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ),
    .Y(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2  (.A1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ),
    .A2(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ),
    .Y(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_b[20] ),
    .B(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__o22a_4 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net182),
    .X(\m_blake2.m_hash256.g_b[20] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X  (.A(net351),
    .B(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(net257),
    .A2(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net395),
    .C1(net179),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net200),
    .A2(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net192),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][20] ),
    .A1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net384),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[21] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ));
 sky130_fd_sc_hd__o21ai_4 \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net182),
    .A2(\m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[22] ),
    .B(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ),
    .A2(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ),
    .Y(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ),
    .B(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .Y(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net183),
    .X(\m_blake2.m_hash256.g_b[22] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net351),
    .A2_N(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net258),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .A2(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net274),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net351),
    .A2(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net180),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][22] ),
    .A1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net383),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[22] ),
    .B(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][22] ),
    .B(net101),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__or4_2 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][22] ),
    .A2(net85),
    .B1(net133),
    .B2(\m_blake2.m_hash256.m_matrix[3][22] ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][22] ),
    .A2(net109),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][22] ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][22] ),
    .A2(net140),
    .B1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net105),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][22] ),
    .A2(net124),
    .B1(net97),
    .B2(\m_blake2.m_hash256.m_matrix[6][22] ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][22] ),
    .A2(net88),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][22] ),
    .C1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][22] ),
    .A2(net112),
    .B1(net137),
    .B2(\m_blake2.m_hash256.m_matrix[2][22] ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][22] ),
    .A2(net129),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][22] ),
    .C1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][22] ),
    .A2(net116),
    .B1(net121),
    .B2(\m_blake2.m_hash256.m_matrix[15][22] ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[23] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__o21ai_4 \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net182),
    .A2(\m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[24] ),
    .B(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net184),
    .X(\m_blake2.m_hash256.g_b[24] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net255),
    .A2(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net380),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net196),
    .A2(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net188),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net353),
    .A2(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net178),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][24] ),
    .A1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net380),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[24] ),
    .B(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ),
    .Y(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__o32a_4 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net100),
    .B2(\m_blake2.m_hash256.m_matrix[0][24] ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][24] ),
    .A2(net118),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][24] ),
    .C1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][24] ),
    .A2(net90),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][24] ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][24] ),
    .A2(net138),
    .B1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][24] ),
    .A2(net114),
    .B1(net98),
    .B2(\m_blake2.m_hash256.m_matrix[6][24] ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][24] ),
    .A2(net130),
    .B1(net134),
    .B2(\m_blake2.m_hash256.m_matrix[3][24] ),
    .C1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][24] ),
    .A2(net86),
    .B1(net110),
    .B2(\m_blake2.m_hash256.m_matrix[7][24] ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][24] ),
    .A2(net126),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][24] ),
    .C1(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][24] ),
    .A2(net146),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][24] ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[25] ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net181),
    .A2(\m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2  (.A1_N(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N ),
    .A2_N(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .B1(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B2(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][25] ),
    .A2(net103),
    .B1(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][25] ),
    .A2(net146),
    .B1(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][25] ),
    .A2(net126),
    .B1(net134),
    .B2(\m_blake2.m_hash256.m_matrix[3][25] ),
    .C1(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][25] ),
    .A2(net90),
    .B1(net114),
    .B2(\m_blake2.m_hash256.m_matrix[5][25] ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][25] ),
    .A2(net130),
    .B1(net118),
    .B2(\m_blake2.m_hash256.m_matrix[13][25] ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][25] ),
    .A2(net94),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][25] ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][25] ),
    .A2(net110),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][25] ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][25] ),
    .A2(net86),
    .B1(net98),
    .B2(\m_blake2.m_hash256.m_matrix[6][25] ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][25] ),
    .A2(net138),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][25] ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_B1 ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[26] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net181),
    .A2(\m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_X ),
    .Y(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.g_b[27] ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net184),
    .A2(\m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B1(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[28] ),
    .B(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_b[28] ),
    .B(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or3b_2_B  (.A(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .C_N(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_A ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net183),
    .X(\m_blake2.m_hash256.g_b[28] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net258),
    .A2(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net381),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net198),
    .A2(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net190),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net353),
    .A2(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net180),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][28] ),
    .A1(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net381),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[29] ),
    .B(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net183),
    .X(\m_blake2.m_hash256.g_b[29] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net360),
    .A2_N(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net257),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o32a_2_X  (.A1(net498),
    .A2(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A3(net274),
    .B1(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net359),
    .A2(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net179),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][29] ),
    .A1(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net397),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[29] ),
    .B(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net177),
    .A2(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net370),
    .X(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net343),
    .A2(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net255),
    .A2(\m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net369),
    .C1(net177),
    .X(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2  (.A1_N(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A1_N ),
    .A2_N(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B2(\m_blake2.m_hash256.g_b[2] ),
    .X(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A2_N_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ),
    .A2(\hash[2]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2_Y ),
    .B1(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A2_N ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[2] ),
    .B(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a22oi_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2  (.A1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1 ),
    .A2(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A2 ),
    .B1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B2(\m_blake2.m_hash256.g_b[30] ),
    .Y(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_Y ));
 sky130_fd_sc_hd__o22a_4 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][30] ),
    .A2(net101),
    .B1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][30] ),
    .A2(net137),
    .B1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net105),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][30] ),
    .A2(net124),
    .B1(net128),
    .B2(\m_blake2.m_hash256.m_matrix[8][30] ),
    .C1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][30] ),
    .A2(net112),
    .B1(net141),
    .B2(\m_blake2.m_hash256.m_matrix[1][30] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][30] ),
    .A2(net96),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][30] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][30] ),
    .A2(net117),
    .B1(net145),
    .B2(\m_blake2.m_hash256.m_matrix[10][30] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][30] ),
    .A2(net109),
    .B1(net88),
    .B2(\m_blake2.m_hash256.m_matrix[14][30] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][30] ),
    .A2(net84),
    .B1(net93),
    .B2(\m_blake2.m_hash256.m_matrix[12][30] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][30] ),
    .A2(net132),
    .B1(net121),
    .B2(\m_blake2.m_hash256.m_matrix[15][30] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net182),
    .X(\m_blake2.m_hash256.g_b[30] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net357),
    .A2_N(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net257),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X  (.A1_N(net192),
    .A2_N(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net274),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net357),
    .A2(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net179),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][30] ),
    .A1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net392),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[30] ),
    .B(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1 ),
    .B(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A2 ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .A2(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X_A ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X  (.A1(net182),
    .A2(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_b[31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][31] ),
    .A1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net396),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X  (.A1(net359),
    .A2(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net396),
    .A2(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B2(net191),
    .C1(net179),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1 ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.g_b[31] ),
    .B(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A ),
    .B(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__o32a_4 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net101),
    .B2(\m_blake2.m_hash256.m_matrix[0][31] ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][31] ),
    .A2(net93),
    .B1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net105),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][31] ),
    .A2(net133),
    .B1(net121),
    .B2(\m_blake2.m_hash256.m_matrix[15][31] ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][31] ),
    .A2(net129),
    .B1(net117),
    .B2(\m_blake2.m_hash256.m_matrix[13][31] ),
    .C1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][31] ),
    .A2(net109),
    .B1(net145),
    .B2(\m_blake2.m_hash256.m_matrix[10][31] ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][31] ),
    .A2(net113),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][31] ),
    .C1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][31] ),
    .A2(net89),
    .B1(net141),
    .B2(\m_blake2.m_hash256.m_matrix[1][31] ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][31] ),
    .A2(net125),
    .B1(net85),
    .B2(\m_blake2.m_hash256.m_matrix[4][31] ),
    .C1(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][31] ),
    .A2(net137),
    .B1(net97),
    .B2(\m_blake2.m_hash256.m_matrix[6][31] ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net178),
    .A2(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net381),
    .X(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net353),
    .A2(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net258),
    .A2(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net381),
    .C1(net180),
    .X(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X ),
    .A2(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_A2 ),
    .B1(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B2(\m_blake2.m_hash256.g_b[3] ),
    .X(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[3] ),
    .B(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[4] ),
    .B(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ba_2_A2  (.A1(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_A ),
    .A2(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1_N(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_C_N ),
    .X(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[4] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net352),
    .A2_N(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net258),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X  (.A1_N(net190),
    .A2_N(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net274),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net352),
    .A2(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net180),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net352),
    .B(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.v_q[4][4] ),
    .A2(net352),
    .B1(net183),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[4] ),
    .B(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[5] ),
    .B(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[5] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net360),
    .A2_N(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net257),
    .X(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X  (.A1_N(net191),
    .A2_N(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ),
    .X(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net359),
    .A2(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net179),
    .X(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net359),
    .B(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.v_q[4][5] ),
    .A2(net359),
    .B1(net182),
    .X(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[5] ),
    .B(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_C_N ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.g_b[6] ),
    .Y(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2  (.A1_N(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X ),
    .A2_N(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .B1(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B2(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_b[6] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net258),
    .A2(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net383),
    .X(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net198),
    .A2(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net190),
    .X(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net351),
    .A2(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net180),
    .X(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net351),
    .B(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.v_q[4][6] ),
    .A2(net351),
    .B1(net183),
    .X(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[7] ),
    .B(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2  (.A1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .A2(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3_2_B  (.A(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .B(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_b[7] ),
    .B(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net182),
    .X(\m_blake2.m_hash256.g_b[7] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X  (.A(net359),
    .B(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(net257),
    .A2(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net396),
    .C1(net179),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net199),
    .A2(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net191),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][7] ),
    .A1(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net396),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_b[8] ),
    .B(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A ),
    .A2(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__nand3_2 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B  (.A(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A ),
    .B(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__and2b_2_B_X ),
    .Y(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_A ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net184),
    .X(\m_blake2.m_hash256.g_b[8] ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(net349),
    .A2_N(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ),
    .B2(net256),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .A2(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net274),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net349),
    .A2(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net178),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][8] ),
    .A1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net376),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.g_b[8] ),
    .B(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__o32ai_4 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y  (.A1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1 ),
    .A2(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2 ),
    .A3(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3 ),
    .B1(net103),
    .B2(\m_blake2.m_hash256.m_matrix[0][8] ),
    .Y(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][8] ),
    .A2(net130),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][8] ),
    .C1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][8] ),
    .A2(net138),
    .B1(net146),
    .B2(\m_blake2.m_hash256.m_matrix[10][8] ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][8] ),
    .A2(net114),
    .B1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][8] ),
    .A2(net110),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][8] ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][8] ),
    .A2(net134),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][8] ),
    .C1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][8] ),
    .A2(net126),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][8] ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][8] ),
    .A2(net118),
    .B1(net98),
    .B2(\m_blake2.m_hash256.m_matrix[6][8] ),
    .C1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][8] ),
    .A2(net86),
    .B1(net90),
    .B2(\m_blake2.m_hash256.m_matrix[14][8] ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_b[9] ),
    .B(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .A2(net104),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.m_matrix[0][9] ),
    .Y(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1 ));
 sky130_fd_sc_hd__nor3_2 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y  (.A(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B ),
    .C(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C ),
    .Y(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][9] ),
    .A2(net118),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][9] ),
    .A2(net130),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][9] ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][9] ),
    .A2(net146),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][9] ),
    .C1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][9] ),
    .A2(net86),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][9] ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][9] ),
    .A2(net114),
    .B1(net98),
    .B2(\m_blake2.m_hash256.m_matrix[6][9] ),
    .C1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][9] ),
    .A2(net90),
    .B1(net138),
    .B2(\m_blake2.m_hash256.m_matrix[2][9] ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][9] ),
    .A2(net110),
    .B1(net134),
    .B2(\m_blake2.m_hash256.m_matrix[3][9] ),
    .C1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][9] ),
    .A2(net126),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][9] ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B  (.A(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ),
    .B(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ),
    .Y(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ),
    .A2(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_C ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_b[9] ),
    .B(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net181),
    .X(\m_blake2.m_hash256.g_b[9] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X  (.A1(net255),
    .A2(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net367),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(net195),
    .A2(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net187),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X  (.A1(net345),
    .A2(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(net177),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[4][9] ),
    .A1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .S(net367),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[0].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[0] ),
    .X(\m_blake2.m_hash256.g_c[0] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[0].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[0] ),
    .X(\m_blake2.m_hash256.g_y[0] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[10].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[10] ),
    .X(\m_blake2.m_hash256.g_c[10] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[10].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[10] ),
    .X(\m_blake2.m_hash256.g_y[10] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[11].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[11] ),
    .X(\m_blake2.m_hash256.g_c[11] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[11].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[11] ),
    .X(\m_blake2.m_hash256.g_y[11] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[12].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[12] ),
    .X(\m_blake2.m_hash256.g_c[12] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[12].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[12] ),
    .X(\m_blake2.m_hash256.g_y[12] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[13].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[13] ),
    .X(\m_blake2.m_hash256.g_c[13] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[13].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[13] ),
    .X(\m_blake2.m_hash256.g_y[13] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[14].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[14] ),
    .X(\m_blake2.m_hash256.g_c[14] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[14].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[14] ),
    .X(\m_blake2.m_hash256.g_y[14] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[15].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[15] ),
    .X(\m_blake2.m_hash256.g_c[15] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[15].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[15] ),
    .X(\m_blake2.m_hash256.g_y[15] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[16].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[16] ),
    .X(\m_blake2.m_hash256.g_c[16] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[16].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[16] ),
    .X(\m_blake2.m_hash256.g_y[16] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[17].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[17] ),
    .X(\m_blake2.m_hash256.g_c[17] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[17].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[17] ),
    .X(\m_blake2.m_hash256.g_y[17] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[18].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[18] ),
    .X(\m_blake2.m_hash256.g_c[18] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[18].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[18] ),
    .X(\m_blake2.m_hash256.g_y[18] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[19].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[19] ),
    .X(\m_blake2.m_hash256.g_c[19] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[19].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[19] ),
    .X(\m_blake2.m_hash256.g_y[19] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[1].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[1] ),
    .X(\m_blake2.m_hash256.g_c[1] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[1].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[1] ),
    .X(\m_blake2.m_hash256.g_y[1] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[20].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[20] ),
    .X(\m_blake2.m_hash256.g_c[20] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[20].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[20] ),
    .X(\m_blake2.m_hash256.g_y[20] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[21].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[21] ),
    .X(\m_blake2.m_hash256.g_c[21] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[21].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[21] ),
    .X(\m_blake2.m_hash256.g_y[21] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[22].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[22] ),
    .X(\m_blake2.m_hash256.g_c[22] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[22].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[22] ),
    .X(\m_blake2.m_hash256.g_y[22] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[23].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[23] ),
    .X(\m_blake2.m_hash256.g_c[23] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[23].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[23] ),
    .X(\m_blake2.m_hash256.g_y[23] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[24].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[24] ),
    .X(\m_blake2.m_hash256.g_c[24] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[24].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[24] ),
    .X(\m_blake2.m_hash256.g_y[24] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[25].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[25] ),
    .X(\m_blake2.m_hash256.g_c[25] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[25].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[25] ),
    .X(\m_blake2.m_hash256.g_y[25] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[26].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[26] ),
    .X(\m_blake2.m_hash256.g_c[26] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[26].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[26] ),
    .X(\m_blake2.m_hash256.g_y[26] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[27].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[27] ),
    .X(\m_blake2.m_hash256.g_c[27] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[27].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[27] ),
    .X(\m_blake2.m_hash256.g_y[27] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[28].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[28] ),
    .X(\m_blake2.m_hash256.g_c[28] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[28].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[28] ),
    .X(\m_blake2.m_hash256.g_y[28] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[29].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[29] ),
    .X(\m_blake2.m_hash256.g_c[29] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[29].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[29] ),
    .X(\m_blake2.m_hash256.g_y[29] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[2].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[2] ),
    .X(\m_blake2.m_hash256.g_c[2] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[2].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[2] ),
    .X(\m_blake2.m_hash256.g_y[2] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[30].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[30] ),
    .X(\m_blake2.m_hash256.g_c[30] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[30].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[30] ),
    .X(\m_blake2.m_hash256.g_y[30] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[31].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[31] ),
    .X(\m_blake2.m_hash256.g_c[31] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[31].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[31] ),
    .X(\m_blake2.m_hash256.g_y[31] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[3].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[3] ),
    .X(\m_blake2.m_hash256.g_c[3] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[3].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[3] ),
    .X(\m_blake2.m_hash256.g_y[3] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[4].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[4] ),
    .X(\m_blake2.m_hash256.g_c[4] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[4].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[4] ),
    .X(\m_blake2.m_hash256.g_y[4] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[5].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[5] ),
    .X(\m_blake2.m_hash256.g_c[5] ));
 sky130_fd_sc_hd__clkbuf_2 \m_blake2.m_hash256.g_buffer[5].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[5] ),
    .X(\m_blake2.m_hash256.g_y[5] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[6].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[6] ),
    .X(\m_blake2.m_hash256.g_c[6] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[6].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[6] ),
    .X(\m_blake2.m_hash256.g_y[6] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[7].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[7] ),
    .X(\m_blake2.m_hash256.g_c[7] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[7].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[7] ),
    .X(\m_blake2.m_hash256.g_y[7] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[8].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[8] ),
    .X(\m_blake2.m_hash256.g_c[8] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[8].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[8] ),
    .X(\m_blake2.m_hash256.g_y[8] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[9].m_c_buf  (.A(\m_blake2.m_hash256.g_c_buf[9] ),
    .X(\m_blake2.m_hash256.g_c[9] ));
 sky130_fd_sc_hd__clkbuf_1 \m_blake2.m_hash256.g_buffer[9].m_y_buf  (.A(\m_blake2.m_hash256.g_y_buf[9] ),
    .X(\m_blake2.m_hash256.g_y[9] ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[0] ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_c_buf[10]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.v_q[8][10] ),
    .A2(net175),
    .B1(\m_blake2.m_hash256.g_c_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net254),
    .X(\m_blake2.m_hash256.g_c_buf[10] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_c_buf[11]_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][11] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B2(\m_blake2.m_hash256.v_q[11][11] ),
    .C1(\m_blake2.m_hash256.g_c_buf[11]_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[11] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_c_buf[11]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net253),
    .Y(\m_blake2.m_hash256.g_c_buf[11]_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][12] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[12] ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net175),
    .B2(\m_blake2.m_hash256.v_q[8][13] ),
    .X(\m_blake2.m_hash256.g_c_buf[13] ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_c_buf[14]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.v_q[8][14] ),
    .A2(net175),
    .B1(\m_blake2.m_hash256.g_c_buf[14]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net253),
    .X(\m_blake2.m_hash256.g_c_buf[14] ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net175),
    .B2(\m_blake2.m_hash256.v_q[8][15] ),
    .X(\m_blake2.m_hash256.g_c_buf[15] ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_c_buf[16]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.v_q[8][16] ),
    .A2(net175),
    .B1(\m_blake2.m_hash256.g_c_buf[16]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net254),
    .X(\m_blake2.m_hash256.g_c_buf[16] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][17] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(\m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_D1 ),
    .X(\m_blake2.m_hash256.g_c_buf[17] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][18] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(\m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_D1 ),
    .X(\m_blake2.m_hash256.g_c_buf[18] ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_c_buf[19]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.v_q[8][19] ),
    .A2(net175),
    .B1(\m_blake2.m_hash256.g_c_buf[19]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net254),
    .X(\m_blake2.m_hash256.g_c_buf[19] ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.v_q[8][1] ),
    .A2(net175),
    .B1(\m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_c_buf[1] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_c_buf[20]_sky130_fd_sc_hd__and2_2_X  (.A(net354),
    .B(\m_blake2.m_hash256.g_c_buf[20]_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_c_buf[20] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][21] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B2(\m_blake2.m_hash256.v_q[11][21] ),
    .C1(\m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[21] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(net169),
    .A2(\m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net251),
    .X(\m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][22] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(\m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_D1 ),
    .X(\m_blake2.m_hash256.g_c_buf[22] ));
 sky130_fd_sc_hd__o311a_1 \m_blake2.m_hash256.g_c_buf[23]_sky130_fd_sc_hd__o311a_2_X  (.A1(net477),
    .A2(\m_blake2.m_hash256.v_q[8][23] ),
    .A3(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .B1(\m_blake2.m_hash256.g_c_buf[23]_sky130_fd_sc_hd__o311a_2_X_B1 ),
    .C1(net355),
    .X(\m_blake2.m_hash256.g_c_buf[23] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][24] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ),
    .B2(\m_blake2.m_hash256.v_q[10][24] ),
    .C1(\m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[24] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(net252),
    .A2(\m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net171),
    .X(\m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.v_q[11][25] ),
    .A2(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_c_buf[25] ));
 sky130_fd_sc_hd__and3_4 \m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X  (.A(net477),
    .B(net355),
    .C(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][26] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[26] ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_c_buf[27]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.v_q[8][27] ),
    .A2(\m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B ),
    .B1(\m_blake2.m_hash256.g_c_buf[27]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_c_buf[27]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_c_buf[27] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][28] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B2(\m_blake2.m_hash256.v_q[11][28] ),
    .C1(\m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[28] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(net170),
    .A2(\m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net251),
    .X(\m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(\m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B ),
    .B2(\m_blake2.m_hash256.v_q[8][29] ),
    .X(\m_blake2.m_hash256.g_c_buf[29] ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[2] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X  (.A1(net355),
    .A2(\m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net253),
    .X(\m_blake2.m_hash256.g_c_buf[30] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][31] ),
    .A2(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ),
    .B1(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ),
    .B2(\m_blake2.m_hash256.v_q[10][31] ),
    .C1(\m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[31] ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(net252),
    .A2(\m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net172),
    .X(\m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_c_buf[3] ));
 sky130_fd_sc_hd__nor2_8 \m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nor2_2_Y  (.A(net388),
    .B(net253),
    .Y(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][4] ),
    .A2(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[4] ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net175),
    .B2(\m_blake2.m_hash256.v_q[8][5] ),
    .X(\m_blake2.m_hash256.g_c_buf[5] ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[6] ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_c_buf[7] ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[8][8] ),
    .A2(net174),
    .B1(\m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_c_buf[8] ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_c_buf[9]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.v_q[8][9] ),
    .A2(net175),
    .B1(\m_blake2.m_hash256.g_c_buf[9]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(net254),
    .X(\m_blake2.m_hash256.g_c_buf[9] ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X  (.A(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_A ),
    .B(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_B ),
    .C(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C ),
    .X(\m_blake2.m_hash256.g_d[0] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[14][0] ),
    .A2(net374),
    .B1(net185),
    .X(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_A ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[15][0] ),
    .A2(net374),
    .B1(net193),
    .X(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(net237),
    .A2(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(net270),
    .B2(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[10] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net237),
    .A2(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net193),
    .A2(\m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net176),
    .C1(net270),
    .X(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net952),
    .A2(net304),
    .B1(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .A2(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[11] ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.v_q[14][11] ),
    .A2(net377),
    .B1(net185),
    .Y(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A1 ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ),
    .A2(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net1140),
    .A2(net305),
    .B1(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net273),
    .A2(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[12] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[6] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[12] ),
    .C1(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net238),
    .A2(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_d[13] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.v_q[13][13] ),
    .A2(net394),
    .B1(net238),
    .C1(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[15][13] ),
    .A2(net275),
    .B1(net176),
    .B2(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2 ),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[12][13] ),
    .A2(net358),
    .B1(net269),
    .C1(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net273),
    .A2(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[14] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[8] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[14] ),
    .C1(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X  (.A(net269),
    .B(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ),
    .C(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ),
    .D(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ),
    .X(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[15] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[9] ),
    .A2(net261),
    .B1(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net238),
    .A2(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net193),
    .A2(\m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net186),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_d[16] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.v_q[13][16] ),
    .A2(net376),
    .B1(net237),
    .C1(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[15][16] ),
    .A2(net275),
    .B1(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net185),
    .C1(net271),
    .X(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[12][16] ),
    .A2(net349),
    .B1(net268),
    .C1(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net270),
    .A2(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[17] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[11] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[17] ),
    .C1(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net237),
    .A2(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X  (.A1_N(net270),
    .A2_N(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_A2_N ),
    .B1(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_d[18] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[15][18] ),
    .A2(net275),
    .B1(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net237),
    .C1(net270),
    .X(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1 ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B2_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[14][18] ),
    .A2(net374),
    .B1(net176),
    .X(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net271),
    .A2(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[19] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[13] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[19] ),
    .C1(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net237),
    .A2(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X  (.A1(net1295),
    .A2(net275),
    .B1(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[1] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[14][1] ),
    .A2(net370),
    .B1(net185),
    .X(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(net237),
    .A2(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net270),
    .X(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[20] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net238),
    .A2(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[14] ),
    .A2(net263),
    .B1(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[21] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net238),
    .A2(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net193),
    .A2(\m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net176),
    .C1(net273),
    .X(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_config.ll_q[21] ),
    .A2(net306),
    .B1(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[22] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_config.ll_q[22] ),
    .A2(net307),
    .B1(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net238),
    .A2(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net194),
    .A2(\m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net176),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[23] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_config.ll_q[23] ),
    .A2(net306),
    .B1(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net239),
    .A2(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net194),
    .A2(\m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net186),
    .C1(net273),
    .X(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net271),
    .A2(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[24] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[18] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ),
    .B2(\m_io.m_config.ll_q[24] ),
    .C1(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ),
    .B(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ),
    .C(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ),
    .D(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ),
    .X(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .A2(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[25] ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.v_q[14][25] ),
    .A2(net368),
    .B1(net185),
    .Y(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A1 ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ),
    .A2(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[19] ),
    .A2(net259),
    .B1(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[26] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net237),
    .A2(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[20] ),
    .A2(net260),
    .B1(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .A2(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[27] ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.v_q[14][27] ),
    .A2(net375),
    .B1(net185),
    .Y(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A1 ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ),
    .A2(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_config.ll_q[27] ),
    .A2(net305),
    .B1(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net273),
    .A2(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[28] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[22] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[28] ),
    .C1(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X  (.A(net269),
    .B(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ),
    .C(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ),
    .D(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ),
    .X(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[29] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net239),
    .A2(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_config.ll_q[29] ),
    .A2(net306),
    .B1(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X  (.A1(net1218),
    .A2(net275),
    .B1(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1 ),
    .X(\m_blake2.m_hash256.g_d[2] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[14][2] ),
    .A2(net369),
    .B1(net176),
    .X(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.v_q[13][2] ),
    .A2(net369),
    .B1(net237),
    .C1(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__o211a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.v_q[12][2] ),
    .A2(net370),
    .B1(net240),
    .B2(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__o221a_2_X_B2 ),
    .C1(net270),
    .X(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net272),
    .A2(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[30] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[24] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ),
    .B2(\m_io.m_config.ll_q[30] ),
    .C1(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net238),
    .A2(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net194),
    .A2(\m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net176),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_d[31] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.v_q[13][31] ),
    .A2(net393),
    .B1(net239),
    .C1(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[15][31] ),
    .A2(net275),
    .B1(net176),
    .B2(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2 ),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[12][31] ),
    .A2(net357),
    .B1(net269),
    .C1(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_d[3] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.v_q[12][3] ),
    .A2(net381),
    .B1(net240),
    .B2(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X_B2 ),
    .C1(net271),
    .X(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[15][3] ),
    .A2(net381),
    .B1(net193),
    .X(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.v_q[13][3] ),
    .A2(net381),
    .B1(net239),
    .C1(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__o211a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[14][3] ),
    .A2(net381),
    .B1(net185),
    .X(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X  (.A(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_A ),
    .B(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_B ),
    .C(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C ),
    .X(\m_blake2.m_hash256.g_d[4] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[14][4] ),
    .A2(net383),
    .B1(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_A ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[15][4] ),
    .A2(net384),
    .B1(net194),
    .X(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(net239),
    .A2(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net273),
    .X(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[15][5] ),
    .A2(net276),
    .B1(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[5] ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.v_q[14][5] ),
    .A2(net394),
    .B1(net186),
    .X(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(net238),
    .A2(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1 ),
    .B2(net273),
    .X(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net273),
    .A2(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[6] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[0] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[6] ),
    .C1(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net1170),
    .A2(net276),
    .B1(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net238),
    .A2(\m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__a221o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ),
    .C1(net273),
    .X(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2 ),
    .B1(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_blake2.m_hash256.g_d[7] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.v_q[13][7] ),
    .A2(net393),
    .B1(net238),
    .C1(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.v_q[15][7] ),
    .A2(net276),
    .B1(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ),
    .B2(net186),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.v_q[12][7] ),
    .A2(net357),
    .B1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ),
    .C1(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_d[8] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(net193),
    .A2(\m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net185),
    .C1(net271),
    .X(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net890),
    .A2(net304),
    .B1(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net270),
    .A2(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[9] ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[3] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[9] ),
    .C1(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net237),
    .A2(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.g_idx_next[0] ),
    .C(net481),
    .X(\m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(net474),
    .Q(\m_blake2.m_hash256.g_idx_next[0] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_idx_next[1] ),
    .B(\m_blake2.m_hash256.g_idx_next[0] ),
    .X(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.g_idx_next[1] ),
    .B(\m_blake2.m_hash256.g_idx_next[0] ),
    .C(net481),
    .X(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__and3b_2 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C  (.A_N(\m_blake2.m_hash256.g_idx_next[0] ),
    .B(net481),
    .C(\m_blake2.m_hash256.g_idx_next[1] ),
    .X(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(net471),
    .Q(\m_blake2.m_hash256.g_idx_next[1] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.g_idx_next[1] ),
    .Y(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.g_idx_next[1] ),
    .A2(\m_blake2.m_hash256.g_idx_next[0] ),
    .B1(\m_blake2.m_hash256.g_idx_next[2] ),
    .X(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1  (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .Y(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__o21ba_2 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N  (.A1(net418),
    .A2(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1_N(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ));
 sky130_fd_sc_hd__or3b_4 \m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A  (.A(\m_blake2.m_hash256.g_idx_next[1] ),
    .B(\m_blake2.m_hash256.g_idx_next[0] ),
    .C_N(net481),
    .X(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1  (.A1(\m_blake2.m_hash256.g_idx_next[2] ),
    .A2(net481),
    .B1_N(net409),
    .X(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X ));
 sky130_fd_sc_hd__and2b_4 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X ),
    .X(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X ),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N  (.A1(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.g_idx_next[0] ),
    .B1_N(\m_blake2.m_hash256.g_idx_next[2] ),
    .X(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__o21ai_4 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1  (.A1(net418),
    .A2(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_1  (.A1(net413),
    .A2(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_1_Y ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.g_idx_next[2] ),
    .B(net481),
    .X(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(net413),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1  (.A(net301),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.g_idx_next[2] ),
    .X(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1  (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(net467),
    .Q(\m_blake2.m_hash256.g_idx_next[2] ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.g_idx_next[2] ),
    .A2(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.g_idx_next[0] ),
    .B1(\m_blake2.m_hash256.g_idx_next[2] ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(net301),
    .A2(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_1  (.A1(net418),
    .A2(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.g_idx_q[0] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(net474),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B  (.A(net444),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand2_2_B  (.A(net445),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ),
    .Y(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net474),
    .A2(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ),
    .B1(net481),
    .Y(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__inv_2_A  (.A(net474),
    .Y(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.g_idx_q[1] ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net469),
    .A2(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net469),
    .A2(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1(net481),
    .Y(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A  (.A(net472),
    .B(net476),
    .Y(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1  (.A(net472),
    .B(net407),
    .Y(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.g_idx_q[2] ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net481),
    .B(net152),
    .C(\m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C ),
    .X(\m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__a21o_2_X  (.A1(net284),
    .A2(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ),
    .B1(net466),
    .X(\m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net18),
    .B2(\m_blake2.m_hash256.m_matrix[0][0] ),
    .X(\m_blake2.m_hash256.g_y_buf[0] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][0] ),
    .A2(net66),
    .B1(net42),
    .B2(\m_blake2.m_hash256.m_matrix[14][0] ),
    .C1(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][0] ),
    .A2(net62),
    .B1(net30),
    .B2(\m_blake2.m_hash256.m_matrix[13][0] ),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][0] ),
    .A2(net78),
    .B1(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][0] ),
    .A2(net26),
    .B1(net54),
    .B2(\m_blake2.m_hash256.m_matrix[10][0] ),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][0] ),
    .A2(net58),
    .B1(net34),
    .B2(\m_blake2.m_hash256.m_matrix[9][0] ),
    .C1(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][0] ),
    .A2(net82),
    .B1(net70),
    .B2(\m_blake2.m_hash256.m_matrix[7][0] ),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][0] ),
    .A2(net50),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][0] ),
    .C1(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][0] ),
    .A2(net38),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][0] ),
    .X(\m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][10] ),
    .A2(net18),
    .B1(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_y_buf[10] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][10] ),
    .A2(net35),
    .B1(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][10] ),
    .A2(net63),
    .B1(net83),
    .B2(\m_blake2.m_hash256.m_matrix[12][10] ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][10] ),
    .A2(net59),
    .B1(net67),
    .B2(\m_blake2.m_hash256.m_matrix[11][10] ),
    .C1(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][10] ),
    .A2(net31),
    .B1(net71),
    .B2(\m_blake2.m_hash256.m_matrix[7][10] ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][10] ),
    .A2(net51),
    .B1(net75),
    .B2(\m_blake2.m_hash256.m_matrix[4][10] ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][10] ),
    .A2(net26),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][10] ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][10] ),
    .A2(net55),
    .B1(net42),
    .B2(\m_blake2.m_hash256.m_matrix[14][10] ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][10] ),
    .A2(net39),
    .B1(net47),
    .B2(\m_blake2.m_hash256.m_matrix[2][10] ),
    .X(\m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net19),
    .B2(\m_blake2.m_hash256.m_matrix[0][11] ),
    .X(\m_blake2.m_hash256.g_y_buf[11] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][11] ),
    .A2(net77),
    .B1(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][11] ),
    .A2(net30),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][11] ),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][11] ),
    .A2(net25),
    .B1(net51),
    .B2(\m_blake2.m_hash256.m_matrix[6][11] ),
    .C1(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][11] ),
    .A2(net61),
    .B1(net39),
    .B2(\m_blake2.m_hash256.m_matrix[5][11] ),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][11] ),
    .A2(net64),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][11] ),
    .C1(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][11] ),
    .A2(net56),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][11] ),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][11] ),
    .A2(net83),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][11] ),
    .C1(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][11] ),
    .A2(net54),
    .B1(net34),
    .B2(\m_blake2.m_hash256.m_matrix[9][11] ),
    .X(\m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][12] ),
    .X(\m_blake2.m_hash256.g_y_buf[12] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][12] ),
    .A2(net56),
    .B1(net28),
    .B2(\m_blake2.m_hash256.m_matrix[13][12] ),
    .C1(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][12] ),
    .A2(net52),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][12] ),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][12] ),
    .A2(net48),
    .B1(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][12] ),
    .A2(net44),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][12] ),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][12] ),
    .A2(net60),
    .B1(net80),
    .B2(\m_blake2.m_hash256.m_matrix[12][12] ),
    .C1(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][12] ),
    .A2(net32),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][12] ),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][12] ),
    .A2(net64),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][12] ),
    .C1(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][12] ),
    .A2(net24),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][12] ),
    .X(\m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][13] ),
    .X(\m_blake2.m_hash256.g_y_buf[13] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][13] ),
    .A2(net48),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][13] ),
    .C1(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][13] ),
    .A2(net60),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][13] ),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][13] ),
    .A2(net28),
    .B1(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][13] ),
    .A2(net32),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][13] ),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][13] ),
    .A2(net36),
    .B1(net44),
    .B2(\m_blake2.m_hash256.m_matrix[2][13] ),
    .C1(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][13] ),
    .A2(net24),
    .B1(net52),
    .B2(\m_blake2.m_hash256.m_matrix[10][13] ),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][13] ),
    .A2(net80),
    .B1(net64),
    .B2(\m_blake2.m_hash256.m_matrix[11][13] ),
    .C1(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][13] ),
    .A2(net56),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][13] ),
    .X(\m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][14] ),
    .X(\m_blake2.m_hash256.g_y_buf[14] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][14] ),
    .A2(net25),
    .B1(net29),
    .B2(\m_blake2.m_hash256.m_matrix[13][14] ),
    .C1(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][14] ),
    .A2(net57),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][14] ),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][14] ),
    .A2(net73),
    .B1(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][14] ),
    .A2(net32),
    .B1(net44),
    .B2(\m_blake2.m_hash256.m_matrix[2][14] ),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][14] ),
    .A2(net61),
    .B1(net52),
    .B2(\m_blake2.m_hash256.m_matrix[10][14] ),
    .C1(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][14] ),
    .A2(net48),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][14] ),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][14] ),
    .A2(net41),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][14] ),
    .C1(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][14] ),
    .A2(net80),
    .B1(net64),
    .B2(\m_blake2.m_hash256.m_matrix[11][14] ),
    .X(\m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][15] ),
    .A2(net17),
    .B1(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_y_buf[15] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][15] ),
    .A2(net25),
    .B1(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][15] ),
    .A2(net49),
    .B1(net45),
    .B2(\m_blake2.m_hash256.m_matrix[2][15] ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][15] ),
    .A2(net29),
    .B1(net37),
    .B2(\m_blake2.m_hash256.m_matrix[5][15] ),
    .C1(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][15] ),
    .A2(net60),
    .B1(net73),
    .B2(\m_blake2.m_hash256.m_matrix[4][15] ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][15] ),
    .A2(net57),
    .B1(net69),
    .B2(\m_blake2.m_hash256.m_matrix[7][15] ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][15] ),
    .A2(net65),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][15] ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][15] ),
    .A2(net53),
    .B1(net81),
    .B2(\m_blake2.m_hash256.m_matrix[12][15] ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][15] ),
    .A2(net33),
    .B1(net41),
    .B2(\m_blake2.m_hash256.m_matrix[14][15] ),
    .X(\m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net18),
    .B2(\m_blake2.m_hash256.m_matrix[0][16] ),
    .X(\m_blake2.m_hash256.g_y_buf[16] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][16] ),
    .A2(net42),
    .B1(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][16] ),
    .A2(net70),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][16] ),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][16] ),
    .A2(net50),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][16] ),
    .C1(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][16] ),
    .A2(net30),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][16] ),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][16] ),
    .A2(net26),
    .B1(net82),
    .B2(\m_blake2.m_hash256.m_matrix[12][16] ),
    .C1(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][16] ),
    .A2(net34),
    .B1(net66),
    .B2(\m_blake2.m_hash256.m_matrix[11][16] ),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][16] ),
    .A2(net58),
    .B1(net54),
    .B2(\m_blake2.m_hash256.m_matrix[10][16] ),
    .C1(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][16] ),
    .A2(net62),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][16] ),
    .X(\m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net18),
    .B2(\m_blake2.m_hash256.m_matrix[0][17] ),
    .X(\m_blake2.m_hash256.g_y_buf[17] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][17] ),
    .A2(net26),
    .B1(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][17] ),
    .A2(net50),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][17] ),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][17] ),
    .A2(net34),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][17] ),
    .C1(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][17] ),
    .A2(net30),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][17] ),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][17] ),
    .A2(net54),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][17] ),
    .C1(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][17] ),
    .A2(net62),
    .B1(net42),
    .B2(\m_blake2.m_hash256.m_matrix[14][17] ),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][17] ),
    .A2(net82),
    .B1(net66),
    .B2(\m_blake2.m_hash256.m_matrix[11][17] ),
    .C1(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][17] ),
    .A2(net58),
    .B1(net70),
    .B2(\m_blake2.m_hash256.m_matrix[7][17] ),
    .X(\m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net19),
    .B2(\m_blake2.m_hash256.m_matrix[0][18] ),
    .X(\m_blake2.m_hash256.g_y_buf[18] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][18] ),
    .A2(net75),
    .B1(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net23),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][18] ),
    .A2(net63),
    .B1(net71),
    .B2(\m_blake2.m_hash256.m_matrix[7][18] ),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][18] ),
    .A2(net59),
    .B1(net47),
    .B2(\m_blake2.m_hash256.m_matrix[2][18] ),
    .C1(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][18] ),
    .A2(net51),
    .B1(net39),
    .B2(\m_blake2.m_hash256.m_matrix[5][18] ),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][18] ),
    .A2(net55),
    .B1(net35),
    .B2(\m_blake2.m_hash256.m_matrix[9][18] ),
    .C1(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][18] ),
    .A2(net26),
    .B1(net31),
    .B2(\m_blake2.m_hash256.m_matrix[13][18] ),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][18] ),
    .A2(net43),
    .B1(net79),
    .B2(\m_blake2.m_hash256.m_matrix[8][18] ),
    .C1(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][18] ),
    .A2(net83),
    .B1(net67),
    .B2(\m_blake2.m_hash256.m_matrix[11][18] ),
    .X(\m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][19] ),
    .X(\m_blake2.m_hash256.g_y_buf[19] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][19] ),
    .A2(net55),
    .B1(net82),
    .B2(\m_blake2.m_hash256.m_matrix[12][19] ),
    .C1(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][19] ),
    .A2(net66),
    .B1(net79),
    .B2(\m_blake2.m_hash256.m_matrix[8][19] ),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][19] ),
    .A2(net74),
    .B1(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][19] ),
    .A2(net51),
    .B1(net47),
    .B2(\m_blake2.m_hash256.m_matrix[2][19] ),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][19] ),
    .A2(net24),
    .B1(net28),
    .B2(\m_blake2.m_hash256.m_matrix[13][19] ),
    .C1(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][19] ),
    .A2(net61),
    .B1(net39),
    .B2(\m_blake2.m_hash256.m_matrix[5][19] ),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][19] ),
    .A2(net34),
    .B1(net43),
    .B2(\m_blake2.m_hash256.m_matrix[14][19] ),
    .C1(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][19] ),
    .A2(net59),
    .B1(net71),
    .B2(\m_blake2.m_hash256.m_matrix[7][19] ),
    .X(\m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net18),
    .B2(\m_blake2.m_hash256.m_matrix[0][1] ),
    .X(\m_blake2.m_hash256.g_y_buf[1] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][1] ),
    .A2(net66),
    .B1(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][1] ),
    .A2(net42),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][1] ),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][1] ),
    .A2(net30),
    .B1(net54),
    .B2(\m_blake2.m_hash256.m_matrix[10][1] ),
    .C1(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][1] ),
    .A2(net62),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][1] ),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][1] ),
    .A2(net50),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][1] ),
    .C1(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][1] ),
    .A2(net82),
    .B1(net70),
    .B2(\m_blake2.m_hash256.m_matrix[7][1] ),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][1] ),
    .A2(net58),
    .B1(net26),
    .B2(\m_blake2.m_hash256.m_matrix[1][1] ),
    .C1(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][1] ),
    .A2(net34),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][1] ),
    .X(\m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][20] ),
    .X(\m_blake2.m_hash256.g_y_buf[20] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][20] ),
    .A2(net52),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][20] ),
    .C1(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][20] ),
    .A2(net32),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][20] ),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][20] ),
    .A2(net56),
    .B1(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][20] ),
    .A2(net28),
    .B1(net64),
    .B2(\m_blake2.m_hash256.m_matrix[11][20] ),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][20] ),
    .A2(net80),
    .B1(net44),
    .B2(\m_blake2.m_hash256.m_matrix[2][20] ),
    .C1(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][20] ),
    .A2(net68),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][20] ),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][20] ),
    .A2(net60),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][20] ),
    .C1(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][20] ),
    .A2(net24),
    .B1(net48),
    .B2(\m_blake2.m_hash256.m_matrix[6][20] ),
    .X(\m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][21] ),
    .X(\m_blake2.m_hash256.g_y_buf[21] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][21] ),
    .A2(net48),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][21] ),
    .C1(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][21] ),
    .A2(net60),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][21] ),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][21] ),
    .A2(net28),
    .B1(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][21] ),
    .A2(net32),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][21] ),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][21] ),
    .A2(net36),
    .B1(net44),
    .B2(\m_blake2.m_hash256.m_matrix[2][21] ),
    .C1(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][21] ),
    .A2(net24),
    .B1(net52),
    .B2(\m_blake2.m_hash256.m_matrix[10][21] ),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][21] ),
    .A2(net80),
    .B1(net64),
    .B2(\m_blake2.m_hash256.m_matrix[11][21] ),
    .C1(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][21] ),
    .A2(net56),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][21] ),
    .X(\m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net17),
    .B2(\m_blake2.m_hash256.m_matrix[0][22] ),
    .X(\m_blake2.m_hash256.g_y_buf[22] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][22] ),
    .A2(net52),
    .B1(net32),
    .B2(\m_blake2.m_hash256.m_matrix[9][22] ),
    .C1(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][22] ),
    .A2(net24),
    .B1(net28),
    .B2(\m_blake2.m_hash256.m_matrix[13][22] ),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][22] ),
    .A2(net72),
    .B1(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][22] ),
    .A2(net60),
    .B1(net69),
    .B2(\m_blake2.m_hash256.m_matrix[7][22] ),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][22] ),
    .A2(net56),
    .B1(net44),
    .B2(\m_blake2.m_hash256.m_matrix[2][22] ),
    .C1(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][22] ),
    .A2(net48),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][22] ),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][22] ),
    .A2(net41),
    .B1(net77),
    .B2(\m_blake2.m_hash256.m_matrix[8][22] ),
    .C1(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][22] ),
    .A2(net80),
    .B1(net64),
    .B2(\m_blake2.m_hash256.m_matrix[11][22] ),
    .X(\m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net17),
    .B2(\m_blake2.m_hash256.m_matrix[0][23] ),
    .X(\m_blake2.m_hash256.g_y_buf[23] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][23] ),
    .A2(net73),
    .B1(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][23] ),
    .A2(net49),
    .B1(net45),
    .B2(\m_blake2.m_hash256.m_matrix[2][23] ),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][23] ),
    .A2(net61),
    .B1(net37),
    .B2(\m_blake2.m_hash256.m_matrix[5][23] ),
    .C1(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][23] ),
    .A2(net25),
    .B1(net29),
    .B2(\m_blake2.m_hash256.m_matrix[13][23] ),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][23] ),
    .A2(net53),
    .B1(net81),
    .B2(\m_blake2.m_hash256.m_matrix[12][23] ),
    .C1(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][23] ),
    .A2(net65),
    .B1(net77),
    .B2(\m_blake2.m_hash256.m_matrix[8][23] ),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][23] ),
    .A2(net33),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][23] ),
    .C1(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][23] ),
    .A2(net57),
    .B1(net69),
    .B2(\m_blake2.m_hash256.m_matrix[7][23] ),
    .X(\m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net18),
    .B2(\m_blake2.m_hash256.m_matrix[0][24] ),
    .X(\m_blake2.m_hash256.g_y_buf[24] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][24] ),
    .A2(net82),
    .B1(net42),
    .B2(\m_blake2.m_hash256.m_matrix[14][24] ),
    .C1(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][24] ),
    .A2(net26),
    .B1(net50),
    .B2(\m_blake2.m_hash256.m_matrix[6][24] ),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][24] ),
    .A2(net46),
    .B1(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][24] ),
    .A2(net62),
    .B1(net34),
    .B2(\m_blake2.m_hash256.m_matrix[9][24] ),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][24] ),
    .A2(net58),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][24] ),
    .C1(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][24] ),
    .A2(net70),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][24] ),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][24] ),
    .A2(net30),
    .B1(net54),
    .B2(\m_blake2.m_hash256.m_matrix[10][24] ),
    .C1(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][24] ),
    .A2(net66),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][24] ),
    .X(\m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][25] ),
    .A2(net18),
    .B1(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_y_buf[25] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][25] ),
    .A2(net26),
    .B1(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][25] ),
    .A2(net50),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][25] ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][25] ),
    .A2(net34),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][25] ),
    .C1(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][25] ),
    .A2(net30),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][25] ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][25] ),
    .A2(net54),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][25] ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][25] ),
    .A2(net58),
    .B1(net70),
    .B2(\m_blake2.m_hash256.m_matrix[7][25] ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][25] ),
    .A2(net62),
    .B1(net42),
    .B2(\m_blake2.m_hash256.m_matrix[14][25] ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][25] ),
    .A2(net82),
    .B1(net66),
    .B2(\m_blake2.m_hash256.m_matrix[11][25] ),
    .X(\m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][26] ),
    .A2(net18),
    .B1(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_y_buf[26] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][26] ),
    .A2(net75),
    .B1(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net23),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][26] ),
    .A2(net62),
    .B1(net70),
    .B2(\m_blake2.m_hash256.m_matrix[7][26] ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][26] ),
    .A2(net58),
    .B1(net47),
    .B2(\m_blake2.m_hash256.m_matrix[2][26] ),
    .C1(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][26] ),
    .A2(net50),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][26] ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][26] ),
    .A2(net83),
    .B1(net67),
    .B2(\m_blake2.m_hash256.m_matrix[11][26] ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][26] ),
    .A2(net27),
    .B1(net31),
    .B2(\m_blake2.m_hash256.m_matrix[13][26] ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][26] ),
    .A2(net55),
    .B1(net35),
    .B2(\m_blake2.m_hash256.m_matrix[9][26] ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][26] ),
    .A2(net42),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][26] ),
    .X(\m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net19),
    .B2(\m_blake2.m_hash256.m_matrix[0][27] ),
    .X(\m_blake2.m_hash256.g_y_buf[27] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][27] ),
    .A2(net35),
    .B1(net71),
    .B2(\m_blake2.m_hash256.m_matrix[7][27] ),
    .C1(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][27] ),
    .A2(net51),
    .B1(net55),
    .B2(\m_blake2.m_hash256.m_matrix[10][27] ),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][27] ),
    .A2(net38),
    .B1(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net23),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][27] ),
    .A2(net67),
    .B1(net79),
    .B2(\m_blake2.m_hash256.m_matrix[8][27] ),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][27] ),
    .A2(net30),
    .B1(net75),
    .B2(\m_blake2.m_hash256.m_matrix[4][27] ),
    .C1(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][27] ),
    .A2(net83),
    .B1(net43),
    .B2(\m_blake2.m_hash256.m_matrix[14][27] ),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][27] ),
    .A2(net58),
    .B1(net27),
    .B2(\m_blake2.m_hash256.m_matrix[1][27] ),
    .C1(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][27] ),
    .A2(net63),
    .B1(net47),
    .B2(\m_blake2.m_hash256.m_matrix[2][27] ),
    .X(\m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][28] ),
    .X(\m_blake2.m_hash256.g_y_buf[28] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][28] ),
    .A2(net56),
    .B1(net28),
    .B2(\m_blake2.m_hash256.m_matrix[13][28] ),
    .C1(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][28] ),
    .A2(net52),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][28] ),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][28] ),
    .A2(net48),
    .B1(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][28] ),
    .A2(net44),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][28] ),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][28] ),
    .A2(net60),
    .B1(net80),
    .B2(\m_blake2.m_hash256.m_matrix[12][28] ),
    .C1(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][28] ),
    .A2(net32),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][28] ),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][28] ),
    .A2(net64),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][28] ),
    .C1(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][28] ),
    .A2(net24),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][28] ),
    .X(\m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][29] ),
    .X(\m_blake2.m_hash256.g_y_buf[29] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][29] ),
    .A2(net56),
    .B1(net44),
    .B2(\m_blake2.m_hash256.m_matrix[2][29] ),
    .C1(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][29] ),
    .A2(net60),
    .B1(net52),
    .B2(\m_blake2.m_hash256.m_matrix[10][29] ),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][29] ),
    .A2(net80),
    .B1(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][29] ),
    .A2(net48),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][29] ),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][29] ),
    .A2(net40),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][29] ),
    .C1(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][29] ),
    .A2(net24),
    .B1(net32),
    .B2(\m_blake2.m_hash256.m_matrix[9][29] ),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][29] ),
    .A2(net28),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][29] ),
    .C1(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][29] ),
    .A2(net65),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][29] ),
    .X(\m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][2] ),
    .A2(net19),
    .B1(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_y_buf[2] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][2] ),
    .A2(net27),
    .B1(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][2] ),
    .A2(net31),
    .B1(net39),
    .B2(\m_blake2.m_hash256.m_matrix[5][2] ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][2] ),
    .A2(net59),
    .B1(net75),
    .B2(\m_blake2.m_hash256.m_matrix[4][2] ),
    .C1(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][2] ),
    .A2(net50),
    .B1(net79),
    .B2(\m_blake2.m_hash256.m_matrix[8][2] ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][2] ),
    .A2(net62),
    .B1(net70),
    .B2(\m_blake2.m_hash256.m_matrix[7][2] ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][2] ),
    .A2(net55),
    .B1(net67),
    .B2(\m_blake2.m_hash256.m_matrix[11][2] ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][2] ),
    .A2(net35),
    .B1(net47),
    .B2(\m_blake2.m_hash256.m_matrix[2][2] ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][2] ),
    .A2(net83),
    .B1(net43),
    .B2(\m_blake2.m_hash256.m_matrix[14][2] ),
    .X(\m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net17),
    .B2(\m_blake2.m_hash256.m_matrix[0][30] ),
    .X(\m_blake2.m_hash256.g_y_buf[30] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][30] ),
    .A2(net61),
    .B1(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][30] ),
    .A2(net29),
    .B1(net65),
    .B2(\m_blake2.m_hash256.m_matrix[11][30] ),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][30] ),
    .A2(net33),
    .B1(net41),
    .B2(\m_blake2.m_hash256.m_matrix[14][30] ),
    .C1(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][30] ),
    .A2(net53),
    .B1(net37),
    .B2(\m_blake2.m_hash256.m_matrix[5][30] ),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][30] ),
    .A2(net25),
    .B1(net69),
    .B2(\m_blake2.m_hash256.m_matrix[7][30] ),
    .C1(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][30] ),
    .A2(net77),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][30] ),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][30] ),
    .A2(net57),
    .B1(net81),
    .B2(\m_blake2.m_hash256.m_matrix[12][30] ),
    .C1(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][30] ),
    .A2(net49),
    .B1(net45),
    .B2(\m_blake2.m_hash256.m_matrix[2][30] ),
    .X(\m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][31] ),
    .A2(net17),
    .B1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_y_buf[31] ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][31] ),
    .A2(net33),
    .B1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][31] ),
    .A2(net49),
    .B1(net53),
    .B2(\m_blake2.m_hash256.m_matrix[10][31] ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][31] ),
    .A2(net25),
    .B1(net69),
    .B2(\m_blake2.m_hash256.m_matrix[7][31] ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][31] ),
    .A2(net57),
    .B1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][31] ),
    .A2(net29),
    .B1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][31] ),
    .A2(net65),
    .B1(net77),
    .B2(\m_blake2.m_hash256.m_matrix[8][31] ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][31] ),
    .A2(net41),
    .B1(net37),
    .B2(\m_blake2.m_hash256.m_matrix[5][31] ),
    .C1(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][31] ),
    .A2(net81),
    .B1(net73),
    .B2(\m_blake2.m_hash256.m_matrix[4][31] ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][31] ),
    .A2(net61),
    .B1(net45),
    .B2(\m_blake2.m_hash256.m_matrix[2][31] ),
    .X(\m_blake2.m_hash256.g_y_buf[31]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net19),
    .B2(\m_blake2.m_hash256.m_matrix[0][3] ),
    .X(\m_blake2.m_hash256.g_y_buf[3] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][3] ),
    .A2(net35),
    .B1(net43),
    .B2(\m_blake2.m_hash256.m_matrix[14][3] ),
    .C1(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][3] ),
    .A2(net59),
    .B1(net71),
    .B2(\m_blake2.m_hash256.m_matrix[7][3] ),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][3] ),
    .A2(net54),
    .B1(net82),
    .B2(\m_blake2.m_hash256.m_matrix[12][3] ),
    .C1(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][3] ),
    .A2(net66),
    .B1(net79),
    .B2(\m_blake2.m_hash256.m_matrix[8][3] ),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][3] ),
    .A2(net27),
    .B1(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net23),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][3] ),
    .A2(net51),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][3] ),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][3] ),
    .A2(net63),
    .B1(net75),
    .B2(\m_blake2.m_hash256.m_matrix[4][3] ),
    .C1(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][3] ),
    .A2(net31),
    .B1(net39),
    .B2(\m_blake2.m_hash256.m_matrix[5][3] ),
    .X(\m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net16),
    .B2(\m_blake2.m_hash256.m_matrix[0][4] ),
    .X(\m_blake2.m_hash256.g_y_buf[4] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][4] ),
    .A2(net60),
    .B1(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][4] ),
    .A2(net44),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][4] ),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][4] ),
    .A2(net48),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][4] ),
    .C1(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][4] ),
    .A2(net32),
    .B1(net80),
    .B2(\m_blake2.m_hash256.m_matrix[12][4] ),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][4] ),
    .A2(net52),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][4] ),
    .C1(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][4] ),
    .A2(net56),
    .B1(net28),
    .B2(\m_blake2.m_hash256.m_matrix[13][4] ),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][4] ),
    .A2(net64),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][4] ),
    .C1(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][4] ),
    .A2(net24),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][4] ),
    .X(\m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][5] ),
    .A2(net16),
    .B1(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.g_y_buf[5] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][5] ),
    .A2(net24),
    .B1(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net20),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][5] ),
    .A2(net48),
    .B1(net44),
    .B2(\m_blake2.m_hash256.m_matrix[2][5] ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][5] ),
    .A2(net32),
    .B1(net72),
    .B2(\m_blake2.m_hash256.m_matrix[4][5] ),
    .C1(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][5] ),
    .A2(net28),
    .B1(net36),
    .B2(\m_blake2.m_hash256.m_matrix[5][5] ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][5] ),
    .A2(net52),
    .B1(net76),
    .B2(\m_blake2.m_hash256.m_matrix[8][5] ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][5] ),
    .A2(net56),
    .B1(net68),
    .B2(\m_blake2.m_hash256.m_matrix[7][5] ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][5] ),
    .A2(net60),
    .B1(net40),
    .B2(\m_blake2.m_hash256.m_matrix[14][5] ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][5] ),
    .A2(net80),
    .B1(net64),
    .B2(\m_blake2.m_hash256.m_matrix[11][5] ),
    .X(\m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net17),
    .B2(\m_blake2.m_hash256.m_matrix[0][6] ),
    .X(\m_blake2.m_hash256.g_y_buf[6] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][6] ),
    .A2(net49),
    .B1(net53),
    .B2(\m_blake2.m_hash256.m_matrix[10][6] ),
    .C1(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][6] ),
    .A2(net33),
    .B1(net65),
    .B2(\m_blake2.m_hash256.m_matrix[11][6] ),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][6] ),
    .A2(net57),
    .B1(net25),
    .B2(\m_blake2.m_hash256.m_matrix[1][6] ),
    .C1(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][6] ),
    .A2(net69),
    .B1(net73),
    .B2(\m_blake2.m_hash256.m_matrix[4][6] ),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][6] ),
    .A2(net81),
    .B1(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][6] ),
    .A2(net37),
    .B1(net45),
    .B2(\m_blake2.m_hash256.m_matrix[2][6] ),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][6] ),
    .A2(net29),
    .B1(net77),
    .B2(\m_blake2.m_hash256.m_matrix[8][6] ),
    .C1(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][6] ),
    .A2(net61),
    .B1(net41),
    .B2(\m_blake2.m_hash256.m_matrix[14][6] ),
    .X(\m_blake2.m_hash256.g_y_buf[6]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net17),
    .B2(\m_blake2.m_hash256.m_matrix[0][7] ),
    .X(\m_blake2.m_hash256.g_y_buf[7] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][7] ),
    .A2(net33),
    .B1(net69),
    .B2(\m_blake2.m_hash256.m_matrix[7][7] ),
    .C1(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][7] ),
    .A2(net49),
    .B1(net73),
    .B2(\m_blake2.m_hash256.m_matrix[4][7] ),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][7] ),
    .A2(net53),
    .B1(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net21),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][7] ),
    .A2(net61),
    .B1(net77),
    .B2(\m_blake2.m_hash256.m_matrix[8][7] ),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][7] ),
    .A2(net41),
    .B1(net37),
    .B2(\m_blake2.m_hash256.m_matrix[5][7] ),
    .C1(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][7] ),
    .A2(net29),
    .B1(net65),
    .B2(\m_blake2.m_hash256.m_matrix[11][7] ),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][7] ),
    .A2(net57),
    .B1(net25),
    .B2(\m_blake2.m_hash256.m_matrix[1][7] ),
    .C1(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][7] ),
    .A2(net81),
    .B1(net45),
    .B2(\m_blake2.m_hash256.m_matrix[2][7] ),
    .X(\m_blake2.m_hash256.g_y_buf[7]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net18),
    .B2(\m_blake2.m_hash256.m_matrix[0][8] ),
    .X(\m_blake2.m_hash256.g_y_buf[8] ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][8] ),
    .A2(net58),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][8] ),
    .C1(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][8] ),
    .A2(net26),
    .B1(net54),
    .B2(\m_blake2.m_hash256.m_matrix[10][8] ),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][8] ),
    .A2(net70),
    .B1(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][8] ),
    .A2(net34),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][8] ),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][8] ),
    .A2(net82),
    .B1(net66),
    .B2(\m_blake2.m_hash256.m_matrix[11][8] ),
    .C1(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][8] ),
    .A2(net30),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][8] ),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][8] ),
    .A2(net62),
    .B1(net42),
    .B2(\m_blake2.m_hash256.m_matrix[14][8] ),
    .C1(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][8] ),
    .A2(net50),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][8] ),
    .X(\m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net18),
    .B2(\m_blake2.m_hash256.m_matrix[0][9] ),
    .X(\m_blake2.m_hash256.g_y_buf[9] ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][9] ),
    .A2(net26),
    .B1(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net22),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][9] ),
    .A2(net30),
    .B1(net82),
    .B2(\m_blake2.m_hash256.m_matrix[12][9] ),
    .C1(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[11][9] ),
    .A2(net66),
    .B1(net38),
    .B2(\m_blake2.m_hash256.m_matrix[5][9] ),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][9] ),
    .A2(net34),
    .B1(net78),
    .B2(\m_blake2.m_hash256.m_matrix[8][9] ),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][9] ),
    .A2(net54),
    .B1(net70),
    .B2(\m_blake2.m_hash256.m_matrix[7][9] ),
    .C1(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][9] ),
    .A2(net50),
    .B1(net74),
    .B2(\m_blake2.m_hash256.m_matrix[4][9] ),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][9] ),
    .A2(net58),
    .B1(net46),
    .B2(\m_blake2.m_hash256.m_matrix[2][9] ),
    .C1(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[15][9] ),
    .A2(net62),
    .B1(net42),
    .B2(\m_blake2.m_hash256.m_matrix[14][9] ),
    .X(\m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[100] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[100] ),
    .A1(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net519),
    .X(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net734),
    .S(net326),
    .X(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__nor2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[100] ),
    .Y(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[101] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[101] ),
    .A1(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net518),
    .X(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net792),
    .S(net325),
    .X(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__or2_2_B  (.A(net494),
    .B(\m_blake2.m_hash256.h_flat[101] ),
    .X(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[102] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[102] ),
    .A1(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net776),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__nand2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[102] ),
    .Y(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[103] ),
    .X(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[103] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[103] ),
    .A1(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net696),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[104] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[104] ),
    .A1(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net744),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__nor2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[104] ),
    .Y(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[105] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[105] ),
    .A1(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net925),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__nand2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[105] ),
    .Y(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[106] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[106] ),
    .A1(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net504),
    .X(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net704),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[106] ),
    .X(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3  (.A1(net470),
    .A2(net475),
    .A3(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(net346),
    .X(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[107] ),
    .X(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[107] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[107] ),
    .A1(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net728),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[108] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[108] ),
    .A1(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net519),
    .X(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net887),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__or2_2_B  (.A(net489),
    .B(\m_blake2.m_hash256.h_flat[108] ),
    .X(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[109] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[109] ),
    .A1(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net518),
    .X(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net833),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__or2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[109] ),
    .X(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[10] ),
    .A1(\m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net507),
    .X(\hash[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net712),
    .S(net316),
    .X(\m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[110] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[110] ),
    .A1(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net739),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__nor2_2_B  (.A(net497),
    .B(\m_blake2.m_hash256.h_flat[110] ),
    .Y(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[111] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[111] ),
    .A1(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net801),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__nor2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[111] ),
    .Y(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[112] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[112] ),
    .A1(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1595),
    .S(net310),
    .X(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__or2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[112] ),
    .X(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[113] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[113] ),
    .A1(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net815),
    .S(net310),
    .X(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__nor2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[113] ),
    .Y(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[114] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[114] ),
    .A1(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net504),
    .X(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net741),
    .S(net312),
    .X(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__nor2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[114] ),
    .Y(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[115] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[115] ),
    .A1(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net714),
    .S(net335),
    .X(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[115] ),
    .X(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B  (.A(net434),
    .B(\m_blake2.m_hash256.h_flat[116] ),
    .X(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2  (.A1(net285),
    .A2(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1_N(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ),
    .X(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[116] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[116] ),
    .A1(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net510),
    .X(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net761),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[117] ),
    .X(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[117] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[117] ),
    .A1(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net751),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[118] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[118] ),
    .A1(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net819),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__nor2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[118] ),
    .Y(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[119] ),
    .X(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[119] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[119] ),
    .A1(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net679),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_X ),
    .A1(net778),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2  (.A1(net531),
    .A2(\m_blake2.m_hash256.h_flat[11] ),
    .B1(\m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2_B2 ),
    .X(\hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[120] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[120] ),
    .A1(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(\m_blake2.m_hash256.h_flat[120] ),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__nor2_2_B  (.A(net489),
    .B(\m_blake2.m_hash256.h_flat[120] ),
    .Y(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[121] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[121] ),
    .A1(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net502),
    .X(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net860),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__nand2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[121] ),
    .Y(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[122] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[122] ),
    .A1(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net847),
    .S(net316),
    .X(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B  (.A(net485),
    .B(\m_blake2.m_hash256.h_flat[122] ),
    .X(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3  (.A1(net469),
    .A2(net474),
    .A3(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(net345),
    .X(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[123] ),
    .X(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[123] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[123] ),
    .A1(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net528),
    .X(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net691),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[124] ),
    .X(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2  (.A1(net288),
    .A2(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(net354),
    .Y(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[124] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[124] ),
    .A1(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net510),
    .X(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1078),
    .S(net326),
    .X(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[125] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[125] ),
    .A1(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1898),
    .S(net335),
    .X(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__nor2_2_B  (.A(net500),
    .B(\m_blake2.m_hash256.h_flat[125] ),
    .Y(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[126] ),
    .X(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[126] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[126] ),
    .A1(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net684),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[127] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[127] ),
    .A1(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net823),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__or2_2_B  (.A(net497),
    .B(\m_blake2.m_hash256.h_flat[127] ),
    .X(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[128] ),
    .A2(net320),
    .B1(\m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net512),
    .B(\m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[128] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[128] ),
    .A1(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net511),
    .X(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.h_flat[128] ),
    .B(net487),
    .Y(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[129] ),
    .A2(net317),
    .B1(\m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net508),
    .B(\m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[129] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[129] ),
    .A1(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__nor2_2_B  (.A(net486),
    .B(\m_blake2.m_hash256.h_flat[129] ),
    .Y(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_X ),
    .A1(net765),
    .S(net323),
    .X(\m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2  (.A1(net510),
    .A2(\m_blake2.m_hash256.h_flat[12] ),
    .B1(\m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2_B2 ),
    .X(\hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[130] ),
    .A2(net320),
    .B1(\m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net512),
    .B(\m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[130] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[130] ),
    .A1(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net507),
    .X(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__nor2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[130] ),
    .Y(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[131] ),
    .A2(net330),
    .B1(\m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net520),
    .B(\m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[131] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[131] ),
    .A1(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__nor2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[131] ),
    .Y(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[132] ),
    .A2(net329),
    .B1(\m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net523),
    .B(\m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[132] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[132] ),
    .A1(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net519),
    .X(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__nor2_2_B  (.A(net493),
    .B(\m_blake2.m_hash256.h_flat[132] ),
    .Y(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[133] ),
    .A2(net340),
    .B1(\m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net537),
    .B(\m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[133] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[133] ),
    .A1(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net530),
    .X(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__nor2_2_B  (.A(net499),
    .B(\m_blake2.m_hash256.h_flat[133] ),
    .Y(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[134] ),
    .A2(net328),
    .B1(\m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net522),
    .B(\m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[134] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[134] ),
    .A1(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__nor2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[134] ),
    .Y(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[135] ),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[135] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[135] ),
    .A1(\m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net872),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net448),
    .A2(net479),
    .A3(\m_blake2.m_hash256.h_flat[136] ),
    .B1(net512),
    .X(\m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[136] ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[136] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net843),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net446),
    .A2(net478),
    .A3(\m_blake2.m_hash256.h_flat[137] ),
    .B1(net507),
    .X(\m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[137] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net767),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__or2_2_B  (.A(net486),
    .B(\m_blake2.m_hash256.h_flat[137] ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net446),
    .A2(net479),
    .A3(\m_blake2.m_hash256.h_flat[138] ),
    .B1(net512),
    .X(\m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[138] ),
    .X(\m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[138] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net742),
    .S(net320),
    .X(\m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net447),
    .A2(net480),
    .A3(\m_blake2.m_hash256.h_flat[139] ),
    .B1(net520),
    .X(\m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__and2_2_B  (.A(net433),
    .B(\m_blake2.m_hash256.h_flat[139] ),
    .X(\m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[139] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net837),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net842),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2  (.A1(net517),
    .A2(\m_blake2.m_hash256.h_flat[13] ),
    .B1(\m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2_B2 ),
    .X(\hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net447),
    .A2(net480),
    .A3(\m_blake2.m_hash256.h_flat[140] ),
    .B1(net522),
    .X(\m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[140] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net762),
    .S(net329),
    .X(\m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[140] ),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net447),
    .A2(net480),
    .A3(\m_blake2.m_hash256.h_flat[141] ),
    .B1(net535),
    .X(\m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__and2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[141] ),
    .X(\m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[141] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net785),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net447),
    .A2(net480),
    .A3(\m_blake2.m_hash256.h_flat[142] ),
    .B1(net522),
    .X(\m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[142] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net806),
    .S(net327),
    .X(\m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[142] ),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[143] ),
    .X(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[143] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[143] ),
    .A1(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net665),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__and2_2_B  (.A(net433),
    .B(\m_blake2.m_hash256.h_flat[144] ),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[144] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[144] ),
    .A1(\m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1267),
    .S(net327),
    .X(\m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[145] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[145] ),
    .A1(\m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net667),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__or2_2_B  (.A(net485),
    .B(\m_blake2.m_hash256.h_flat[145] ),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[146] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[146] ),
    .A1(\m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net512),
    .X(\m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net700),
    .S(net320),
    .X(\m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__or2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[146] ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[147] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[147] ),
    .A1(\m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net802),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__or2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[147] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[148] ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[148] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[148] ),
    .A1(\m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net523),
    .X(\m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net661),
    .S(net329),
    .X(\m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__and2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[149] ),
    .X(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[149] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[149] ),
    .A1(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net725),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[14] ),
    .A1(\m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net530),
    .X(\hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net713),
    .S(net335),
    .X(\m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__or2_2_B  (.A(net500),
    .B(\m_blake2.m_hash256.h_flat[14] ),
    .X(\m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__and2_2_B  (.A(net436),
    .B(\m_blake2.m_hash256.h_flat[150] ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[150] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[150] ),
    .A1(\m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net520),
    .X(\m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1047),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[151] ),
    .X(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[151] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[151] ),
    .A1(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net662),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[152] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[152] ),
    .A1(\m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net520),
    .X(\m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net705),
    .S(net327),
    .X(\m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[152] ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__and2_2_B  (.A(net430),
    .B(\m_blake2.m_hash256.h_flat[153] ),
    .X(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[153] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[153] ),
    .A1(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net721),
    .S(net317),
    .X(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[154] ),
    .X(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[154] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[154] ),
    .A1(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net512),
    .X(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net671),
    .S(net320),
    .X(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__and2_2_B  (.A(net433),
    .B(\m_blake2.m_hash256.h_flat[155] ),
    .X(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[155] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[155] ),
    .A1(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net735),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[156] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[156] ),
    .A1(\m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net523),
    .X(\m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net698),
    .S(net329),
    .X(\m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__or2_2_B  (.A(net493),
    .B(\m_blake2.m_hash256.h_flat[156] ),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__and2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[157] ),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[157] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[157] ),
    .A1(\m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net719),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[158] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[158] ),
    .A1(\m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net522),
    .X(\m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net717),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__or2_2_B  (.A(net499),
    .B(\m_blake2.m_hash256.h_flat[158] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[159] ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__mux2_1_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[159] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[159] ),
    .A1(\m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1286),
    .S(net338),
    .X(\m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[15] ),
    .A1(\m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net530),
    .X(\hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net866),
    .S(net335),
    .X(\m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__or2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[15] ),
    .X(\m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[160] ),
    .X(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[160] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[160] ),
    .A1(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net520),
    .X(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1696),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__and2_2_B  (.A(net431),
    .B(\m_blake2.m_hash256.h_flat[161] ),
    .X(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[161] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[161] ),
    .A1(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net508),
    .X(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net809),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net654),
    .A2(net319),
    .B1(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[162] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[162] ),
    .A1(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net512),
    .X(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[162] ),
    .X(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net197),
    .A2(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net187),
    .X(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net740),
    .A2(net327),
    .B1(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[163] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[163] ),
    .A1(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__or2_2_B  (.A(net493),
    .B(\m_blake2.m_hash256.h_flat[163] ),
    .X(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__and2_2_B  (.A(net436),
    .B(\m_blake2.m_hash256.h_flat[164] ),
    .X(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[164] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[164] ),
    .A1(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net523),
    .X(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net688),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__and2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[165] ),
    .X(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[165] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[165] ),
    .A1(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net729),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[166] ),
    .X(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[166] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[166] ),
    .A1(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net531),
    .X(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1021),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net658),
    .A2(net338),
    .B1(\m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net534),
    .B(\m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[167] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[167] ),
    .A1(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net534),
    .X(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__or2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[167] ),
    .X(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[168] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[168] ),
    .A1(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net791),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__nand2_2_B  (.A(net433),
    .B(\m_blake2.m_hash256.h_flat[168] ),
    .Y(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__and2_2_B  (.A(net430),
    .B(\m_blake2.m_hash256.h_flat[169] ),
    .X(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[169] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[169] ),
    .A1(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net737),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__and2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[16] ),
    .X(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net782),
    .S(net310),
    .X(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__o22a_2_A2  (.A1(net501),
    .A2(\m_blake2.m_hash256.h_flat[16] ),
    .B1(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__o22a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__o22a_2_A2_B2 ),
    .X(\m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__and3_2_C  (.A(net448),
    .B(net479),
    .C(\m_blake2.m_hash256.h_flat[170] ),
    .X(\m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net513),
    .X(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[170] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net730),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__nand2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[170] ),
    .Y(\m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__and3_2_C  (.A(net447),
    .B(net480),
    .C(\m_blake2.m_hash256.h_flat[171] ),
    .X(\m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net521),
    .X(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[171] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net780),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[171] ),
    .X(\m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[172] ),
    .X(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[172] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[172] ),
    .A1(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net523),
    .X(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1563),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[173] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[173] ),
    .A1(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net666),
    .S(net340),
    .X(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[173] ),
    .X(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net199),
    .A2(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net192),
    .X(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[174] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[174] ),
    .A1(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net522),
    .X(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net657),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[174] ),
    .X(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net448),
    .A2(net480),
    .A3(\m_blake2.m_hash256.h_flat[175] ),
    .B1(net534),
    .X(\m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[175] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net816),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__nand2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[175] ),
    .Y(\m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[176] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[176] ),
    .A1(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net763),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__or2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[176] ),
    .X(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__and2_2_B  (.A(net430),
    .B(\m_blake2.m_hash256.h_flat[177] ),
    .X(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[177] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[177] ),
    .A1(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net736),
    .S(net316),
    .X(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[178] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[178] ),
    .A1(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net513),
    .X(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net726),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__or2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[178] ),
    .X(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__and2_2_B  (.A(net433),
    .B(\m_blake2.m_hash256.h_flat[179] ),
    .X(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[179] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[179] ),
    .A1(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1250),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__and2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[17] ),
    .X(\m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[17] ),
    .A1(\m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net845),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[180] ),
    .X(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[180] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[180] ),
    .A1(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net531),
    .X(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net899),
    .S(net341),
    .X(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[181] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[181] ),
    .A1(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net759),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__nand2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[181] ),
    .Y(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[182] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[182] ),
    .A1(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net522),
    .X(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net863),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__nand2_2_B  (.A(net436),
    .B(\m_blake2.m_hash256.h_flat[182] ),
    .Y(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[183] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[183] ),
    .A1(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net865),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__nand2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[183] ),
    .Y(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[184] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[184] ),
    .A1(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net664),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[184] ),
    .X(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[185] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[185] ),
    .A1(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net770),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__or2_2_B  (.A(net485),
    .B(\m_blake2.m_hash256.h_flat[185] ),
    .X(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[186] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[186] ),
    .A1(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net512),
    .X(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net827),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__nand2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[186] ),
    .Y(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[187] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[187] ),
    .A1(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net516),
    .X(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net786),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__or2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[187] ),
    .X(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[188] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[188] ),
    .A1(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net532),
    .X(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1824),
    .S(net330),
    .X(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[188] ),
    .X(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[189] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[189] ),
    .A1(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net536),
    .X(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net805),
    .S(net340),
    .X(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__nand2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[189] ),
    .Y(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__and2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[18] ),
    .X(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[18] ),
    .A1(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net504),
    .X(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net727),
    .S(net312),
    .X(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[190] ),
    .X(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[190] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[190] ),
    .A1(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net531),
    .X(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net675),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[191] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[191] ),
    .A1(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net534),
    .X(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net682),
    .S(net338),
    .X(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__or2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[191] ),
    .X(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net908),
    .A2(net321),
    .B1(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[192] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[192] ),
    .A1(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__or2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[192] ),
    .X(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net711),
    .A2(net315),
    .B1(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[193] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[193] ),
    .A1(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__or2_2_B  (.A(net485),
    .B(\m_blake2.m_hash256.h_flat[193] ),
    .X(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__and2_2_B  (.A(net430),
    .B(\m_blake2.m_hash256.h_flat[194] ),
    .X(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[194] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[194] ),
    .A1(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net512),
    .X(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1109),
    .S(net317),
    .X(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net850),
    .A2(net327),
    .B1(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[195] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[195] ),
    .A1(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net516),
    .X(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__or2_2_B  (.A(net493),
    .B(\m_blake2.m_hash256.h_flat[195] ),
    .X(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__and2_2_B  (.A(net436),
    .B(\m_blake2.m_hash256.h_flat[196] ),
    .X(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[196] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[196] ),
    .A1(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net521),
    .X(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net738),
    .S(net329),
    .X(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net652),
    .A2(net339),
    .B1(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[197] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[197] ),
    .A1(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net536),
    .X(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__or2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[197] ),
    .X(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[198] ),
    .X(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[198] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[198] ),
    .A1(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net531),
    .X(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1135),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net653),
    .A2(net337),
    .B1(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[199] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[199] ),
    .A1(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__or2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[199] ),
    .X(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1003),
    .S(net335),
    .X(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2  (.A1(net530),
    .A2(\m_blake2.m_hash256.h_flat[19] ),
    .B1(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_B2 ),
    .X(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[19] ),
    .X(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__and3_2_C  (.A(net448),
    .B(net479),
    .C(\m_blake2.m_hash256.h_flat[200] ),
    .X(\m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[200] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net784),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__or2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[200] ),
    .X(\m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and2_2_B  (.A(net430),
    .B(\m_blake2.m_hash256.h_flat[201] ),
    .X(\m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and3_2_C  (.A(net446),
    .B(net478),
    .C(\m_blake2.m_hash256.h_flat[201] ),
    .X(\m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[201] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net799),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__and2_2_B  (.A(net431),
    .B(\m_blake2.m_hash256.h_flat[202] ),
    .X(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[202] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[202] ),
    .A1(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net508),
    .X(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net677),
    .S(net317),
    .X(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C  (.A(net447),
    .B(net480),
    .C(\m_blake2.m_hash256.h_flat[203] ),
    .X(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net520),
    .X(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[203] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net800),
    .S(net327),
    .X(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[203] ),
    .X(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(net274),
    .A2_N(\m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net255),
    .X(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[204] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[204] ),
    .A1(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net523),
    .X(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(\m_blake2.m_hash256.h_flat[204] ),
    .S(net341),
    .X(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__or2_2_B  (.A(net499),
    .B(\m_blake2.m_hash256.h_flat[204] ),
    .X(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[205] ),
    .X(\m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and3_2_C  (.A(net447),
    .B(net480),
    .C(\m_blake2.m_hash256.h_flat[205] ),
    .X(\m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[205] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net699),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[206] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[206] ),
    .A1(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net522),
    .X(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net826),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[206] ),
    .X(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__and3_2_C  (.A(net447),
    .B(net480),
    .C(\m_blake2.m_hash256.h_flat[207] ),
    .X(\m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net534),
    .X(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[207] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net692),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__or2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[207] ),
    .X(\m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[208] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[208] ),
    .A1(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1104),
    .S(net327),
    .X(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[208] ),
    .X(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[209] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[209] ),
    .A1(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net752),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__or2_2_B  (.A(net485),
    .B(\m_blake2.m_hash256.h_flat[209] ),
    .X(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__and2_2_B  (.A(net434),
    .B(\m_blake2.m_hash256.h_flat[20] ),
    .X(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net796),
    .S(net323),
    .X(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2  (.A1(net510),
    .A2(\m_blake2.m_hash256.h_flat[20] ),
    .B1(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_B2 ),
    .X(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[210] ),
    .X(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[210] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[210] ),
    .A1(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net508),
    .X(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net766),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[211] ),
    .X(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[211] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[211] ),
    .A1(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net521),
    .X(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1086),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[212] ),
    .X(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[212] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[212] ),
    .A1(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net532),
    .X(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net964),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__and2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[213] ),
    .X(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[213] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[213] ),
    .A1(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net764),
    .S(net340),
    .X(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[214] ),
    .X(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[214] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[214] ),
    .A1(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net522),
    .X(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1468),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[215] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[215] ),
    .A1(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net760),
    .S(net338),
    .X(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__or2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[215] ),
    .X(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[216] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[216] ),
    .A1(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net520),
    .X(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net668),
    .S(net327),
    .X(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[216] ),
    .X(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[217] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[217] ),
    .A1(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net747),
    .S(net317),
    .X(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__or2_2_B  (.A(net485),
    .B(\m_blake2.m_hash256.h_flat[217] ),
    .X(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[218] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[218] ),
    .A1(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net513),
    .X(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net697),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__or2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[218] ),
    .X(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[219] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[219] ),
    .A1(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net659),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__or2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[219] ),
    .X(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[21] ),
    .X(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[21] ),
    .A1(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net807),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[220] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[220] ),
    .A1(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net532),
    .X(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1381),
    .S(net329),
    .X(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[220] ),
    .X(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__and2_2_B  (.A(net442),
    .B(\m_blake2.m_hash256.h_flat[221] ),
    .X(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[221] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[221] ),
    .A1(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net536),
    .X(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net841),
    .S(net340),
    .X(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[222] ),
    .X(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[222] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[222] ),
    .A1(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net531),
    .X(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net846),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[223] ),
    .X(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net199),
    .A2(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net257),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[223] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[223] ),
    .A1(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net534),
    .X(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net716),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.h_flat[224] ),
    .A2(net321),
    .B1(\m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net514),
    .B(\m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[224] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[224] ),
    .A1(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net520),
    .X(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__nor2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[224] ),
    .Y(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[225] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[225] ),
    .A1(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net508),
    .X(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net810),
    .S(net317),
    .X(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__nand2_2_B  (.A(net431),
    .B(\m_blake2.m_hash256.h_flat[225] ),
    .Y(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[226] ),
    .X(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[226] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[226] ),
    .A1(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net513),
    .X(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net708),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__a21o_2_A1  (.A1(net680),
    .A2(net327),
    .B1(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[227] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[227] ),
    .A1(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[227] ),
    .X(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net198),
    .A2(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net190),
    .X(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net804),
    .A2(net329),
    .B1(\m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B2(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__a22o_2_A1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(net523),
    .B(\m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__a22o_2_A1_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[228] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[228] ),
    .A1(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net523),
    .X(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__nor2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[228] ),
    .Y(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[229] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[229] ),
    .A1(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net536),
    .X(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net913),
    .S(net340),
    .X(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__nand2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[229] ),
    .Y(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__and2_2_B  (.A(net442),
    .B(\m_blake2.m_hash256.h_flat[22] ),
    .X(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[22] ),
    .A1(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net530),
    .X(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net694),
    .S(net335),
    .X(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__and2_2_B  (.A(net436),
    .B(\m_blake2.m_hash256.h_flat[230] ),
    .X(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[230] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[230] ),
    .A1(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net531),
    .X(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1556),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[231] ),
    .X(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[231] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[231] ),
    .A1(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net788),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net446),
    .A2(net479),
    .A3(\m_blake2.m_hash256.h_flat[232] ),
    .B1(net514),
    .X(\m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[232] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net885),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__nor2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[232] ),
    .Y(\m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__and2_2_B  (.A(net430),
    .B(\m_blake2.m_hash256.h_flat[233] ),
    .X(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[233] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[233] ),
    .A1(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net508),
    .X(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net722),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[234] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[234] ),
    .A1(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net513),
    .X(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net756),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[234] ),
    .Y(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .A2(\m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net274),
    .X(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C  (.A(net447),
    .B(net480),
    .C(\m_blake2.m_hash256.h_flat[235] ),
    .X(\m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C_X ),
    .A1(\m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net520),
    .X(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[235] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net808),
    .S(net330),
    .X(\m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__nor2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[235] ),
    .Y(\m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net447),
    .A2(\m_blake2.m_hash256.fsm_q[4] ),
    .A3(\m_blake2.m_hash256.h_flat[236] ),
    .B1(net532),
    .X(\m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[236] ),
    .X(\m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[236] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net777),
    .S(net341),
    .X(\m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__and2_2_B  (.A(net439),
    .B(\m_blake2.m_hash256.h_flat[237] ),
    .X(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[237] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[237] ),
    .A1(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net537),
    .X(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net693),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[238] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[238] ),
    .A1(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net522),
    .X(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net754),
    .S(net328),
    .X(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[238] ),
    .X(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[239] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[239] ),
    .A1(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net748),
    .S(net337),
    .X(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[239] ),
    .Y(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .A2(\m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ),
    .X(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[23] ),
    .X(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[23] ),
    .A1(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net530),
    .X(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net718),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__and2_2_B  (.A(net433),
    .B(\m_blake2.m_hash256.h_flat[240] ),
    .X(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[240] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[240] ),
    .A1(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net514),
    .X(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net701),
    .S(net321),
    .X(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__and2_2_B  (.A(net430),
    .B(\m_blake2.m_hash256.h_flat[241] ),
    .X(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[241] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[241] ),
    .A1(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net506),
    .X(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net753),
    .S(net315),
    .X(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__and2_2_B  (.A(net432),
    .B(\m_blake2.m_hash256.h_flat[242] ),
    .X(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[242] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[242] ),
    .A1(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net513),
    .X(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net859),
    .S(net319),
    .X(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__and2_2_B  (.A(net433),
    .B(\m_blake2.m_hash256.h_flat[243] ),
    .X(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[243] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[243] ),
    .A1(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net521),
    .X(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1376),
    .S(net322),
    .X(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__and2_2_B  (.A(net441),
    .B(\m_blake2.m_hash256.h_flat[244] ),
    .X(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[244] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[244] ),
    .A1(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net532),
    .X(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net900),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[245] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[245] ),
    .A1(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net535),
    .X(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net838),
    .S(net339),
    .X(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B  (.A(net499),
    .B(\m_blake2.m_hash256.h_flat[245] ),
    .Y(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .A2(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ),
    .X(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[246] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[246] ),
    .A1(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net522),
    .X(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1657),
    .S(net336),
    .X(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__nor2_2_B  (.A(net499),
    .B(\m_blake2.m_hash256.h_flat[246] ),
    .Y(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[247] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[247] ),
    .A1(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net811),
    .S(net338),
    .X(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B  (.A(net498),
    .B(\m_blake2.m_hash256.h_flat[247] ),
    .Y(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .A2(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ),
    .X(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net758),
    .A2(net327),
    .B1(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__a22o_2_A1_B1 ),
    .B2(net520),
    .X(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[248] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[248] ),
    .A1(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__or2_2_B  (.A(net491),
    .B(\m_blake2.m_hash256.h_flat[248] ),
    .X(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net732),
    .A2(net317),
    .B1(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__a22o_2_A1_B1 ),
    .B2(net508),
    .X(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[249] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[249] ),
    .A1(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net508),
    .X(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B  (.A(net486),
    .B(\m_blake2.m_hash256.h_flat[249] ),
    .X(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net195),
    .A2(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net187),
    .X(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[24] ),
    .A1(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(\m_blake2.m_hash256.h_flat[24] ),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__or2_2_B  (.A(net489),
    .B(\m_blake2.m_hash256.h_flat[24] ),
    .X(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net1072),
    .A2(net319),
    .B1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__a22o_2_A1_B1 ),
    .B2(net512),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[250] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.h_flat[250] ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(net487),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2  (.A1(net487),
    .A2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A3(net274),
    .B1(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_X ));
 sky130_fd_sc_hd__nand2_8 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__inv_6 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__inv_2_Y  (.A(net469),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__nor2_8 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(net407),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y  (.A(net467),
    .B(net476),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B ),
    .B(net249),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B  (.A(net471),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(net475),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B  (.A(net344),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ),
    .C(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__nand2_8 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand2_2_B  (.A(net471),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B  (.A(net473),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__o211a_2_C1  (.A1(net449),
    .A2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .C1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__o211a_2_C1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__or2_4 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1  (.A(net473),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B  (.A(net304),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__xor2_2_X  (.A(net467),
    .B(net475),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[250] ),
    .A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net513),
    .X(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net669),
    .A2(net322),
    .B1(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__a22o_2_A1_B1 ),
    .B2(net515),
    .X(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[251] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[251] ),
    .A1(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net515),
    .X(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B  (.A(net488),
    .B(\m_blake2.m_hash256.h_flat[251] ),
    .X(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net196),
    .A2(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net189),
    .X(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net1856),
    .A2(net329),
    .B1(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__a22o_2_A1_B1 ),
    .B2(net521),
    .X(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[252] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[252] ),
    .A1(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net532),
    .X(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__or2_2_B  (.A(net492),
    .B(\m_blake2.m_hash256.h_flat[252] ),
    .X(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net1348),
    .A2(net339),
    .B1(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__a22o_2_A1_B1 ),
    .B2(net535),
    .X(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[253] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.h_flat[253] ),
    .Y(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(net499),
    .B(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[253] ),
    .A1(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net536),
    .X(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__a22o_2_A1  (.A1(net774),
    .A2(net336),
    .B1(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__a22o_2_A1_B1 ),
    .B2(net531),
    .X(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[254] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[254] ),
    .A1(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net531),
    .X(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__nor2_2_B  (.A(net499),
    .B(\m_blake2.m_hash256.h_flat[254] ),
    .Y(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__a32o_2_B1  (.A1(net534),
    .A2(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__a32o_2_B1_A2 ),
    .A3(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__a32o_2_B1_A3 ),
    .B1(net645),
    .B2(net338),
    .X(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[255] ),
    .X(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[255] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[255] ),
    .A1(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net533),
    .X(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[25] ),
    .A1(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net502),
    .X(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1499),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__or2_2_B  (.A(net486),
    .B(\m_blake2.m_hash256.h_flat[25] ),
    .X(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__and2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[26] ),
    .X(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[26] ),
    .A1(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net504),
    .X(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net768),
    .S(net312),
    .X(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[27] ),
    .A1(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net530),
    .X(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net687),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[27] ),
    .X(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[28] ),
    .X(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[28] ),
    .A1(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net510),
    .X(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1235),
    .S(net326),
    .X(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[29] ),
    .A1(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1017),
    .S(net325),
    .X(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__or2_2_B  (.A(net494),
    .B(\m_blake2.m_hash256.h_flat[29] ),
    .X(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[30] ),
    .A1(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net530),
    .X(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net835),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__or2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[30] ),
    .X(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[31] ),
    .X(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[31] ),
    .A1(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net529),
    .X(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net683),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[32] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[32] ),
    .A1(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net511),
    .X(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1445),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B  (.A(net486),
    .B(\m_blake2.m_hash256.h_flat[32] ),
    .X(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2  (.A1(net290),
    .A2(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net278),
    .C1(\hash[0]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ),
    .X(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[33] ),
    .X(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net289),
    .A2(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ),
    .X(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[33] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[33] ),
    .A1(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net686),
    .S(net312),
    .X(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[34] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[34] ),
    .A1(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net504),
    .X(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net775),
    .S(net312),
    .X(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[34] ),
    .Y(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1  (.A1(net266),
    .A2(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net267),
    .X(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__nand2_4 \m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(net475),
    .Y(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B  (.A(net440),
    .B(\m_blake2.m_hash256.h_flat[35] ),
    .X(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net293),
    .A2(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ),
    .X(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[35] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[35] ),
    .A1(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net529),
    .X(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net672),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[36] ),
    .X(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2  (.A1(net295),
    .A2(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(net350),
    .Y(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[36] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[36] ),
    .A1(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net519),
    .X(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net690),
    .S(net326),
    .X(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B  (.A(net435),
    .B(\m_blake2.m_hash256.h_flat[37] ),
    .X(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net295),
    .A2(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .X(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[37] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[37] ),
    .A1(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net518),
    .X(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net707),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[38] ),
    .X(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net292),
    .A2(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ),
    .C1(net356),
    .X(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[38] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[38] ),
    .A1(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net720),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[39] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[39] ),
    .A1(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net529),
    .X(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net723),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[39] ),
    .X(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net286),
    .A2(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net293),
    .X(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[40] ),
    .X(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21boi_1 \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2  (.A1(net290),
    .A2(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1_N(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_X ),
    .Y(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[40] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[40] ),
    .A1(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net673),
    .S(net314),
    .X(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[41] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[41] ),
    .A1(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net504),
    .X(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net825),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[41] ),
    .Y(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1  (.A1(net400),
    .A2(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net267),
    .C1(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[42] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[42] ),
    .A1(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net504),
    .X(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net813),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[42] ),
    .X(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net277),
    .A2(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net289),
    .X(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[43] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[43] ),
    .A1(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net529),
    .X(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net822),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[43] ),
    .Y(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net266),
    .C1(net389),
    .X(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B  (.A(net434),
    .B(\m_blake2.m_hash256.h_flat[44] ),
    .X(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net291),
    .A2(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .X(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[44] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[44] ),
    .A1(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net519),
    .X(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1068),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[45] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[45] ),
    .A1(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net518),
    .X(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net745),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[45] ),
    .X(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net295),
    .A2(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net406),
    .X(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[46] ),
    .X(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net292),
    .A2(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ),
    .C1(net356),
    .X(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[46] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[46] ),
    .A1(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net674),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[47] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[47] ),
    .A1(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net529),
    .X(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net832),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[47] ),
    .Y(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o211ai_1 \m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ),
    .C1(net389),
    .Y(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[48] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[48] ),
    .A1(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net509),
    .X(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net893),
    .S(net310),
    .X(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B  (.A(net486),
    .B(\m_blake2.m_hash256.h_flat[48] ),
    .X(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net284),
    .A2(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net289),
    .X(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or3_2_C  (.A(net346),
    .B(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .C(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[49] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[49] ),
    .A1(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net773),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[49] ),
    .Y(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o211ai_1 \m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ),
    .C1(net362),
    .Y(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[50] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[50] ),
    .A1(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net923),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[50] ),
    .Y(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o211ai_1 \m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ),
    .C1(net363),
    .Y(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[51] ),
    .X(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net293),
    .A2(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .C1(net356),
    .X(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[51] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[51] ),
    .A1(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net529),
    .X(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net678),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[52] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[52] ),
    .A1(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net510),
    .X(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net771),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B  (.A(net434),
    .B(\m_blake2.m_hash256.h_flat[52] ),
    .Y(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net266),
    .C1(net372),
    .X(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[53] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[53] ),
    .A1(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net779),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[53] ),
    .X(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net288),
    .A2(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net295),
    .X(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[54] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[54] ),
    .A1(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net702),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[54] ),
    .X(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2  (.A1(net292),
    .A2(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1_N(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ),
    .X(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[55] ),
    .X(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1  (.A1(net286),
    .A2(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net292),
    .C1(net355),
    .X(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[55] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[55] ),
    .A1(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net663),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[56] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[56] ),
    .A1(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(\m_blake2.m_hash256.h_flat[56] ),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B  (.A(net489),
    .B(\m_blake2.m_hash256.h_flat[56] ),
    .Y(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22ai_1 \m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net400),
    .Y(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[57] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[57] ),
    .A1(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net864),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[57] ),
    .Y(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22ai_1 \m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net400),
    .Y(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__and2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[58] ),
    .X(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[58] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[58] ),
    .A1(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net749),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[59] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[59] ),
    .A1(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net528),
    .X(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net733),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[59] ),
    .X(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2  (.A1(net293),
    .A2(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .C1(net356),
    .Y(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[60] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[60] ),
    .A1(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net510),
    .X(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net803),
    .S(net323),
    .X(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__nor2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[60] ),
    .Y(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[61] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[61] ),
    .A1(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net787),
    .S(net325),
    .X(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[61] ),
    .Y(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2  (.A1(net267),
    .A2(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ),
    .C1(net379),
    .X(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[62] ),
    .X(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net292),
    .A2(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .C1(net356),
    .X(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[62] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[62] ),
    .A1(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net685),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[63] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[63] ),
    .A1(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net818),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[63] ),
    .X(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2  (.A1(net293),
    .A2(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .C1(net356),
    .Y(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__and2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[64] ),
    .X(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[64] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[64] ),
    .A1(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net511),
    .X(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1647),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[65] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[65] ),
    .A1(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net772),
    .S(net310),
    .X(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__or2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[65] ),
    .X(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[66] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[66] ),
    .A1(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net812),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__nand2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[66] ),
    .Y(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[67] ),
    .X(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[67] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[67] ),
    .A1(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net676),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[68] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[68] ),
    .A1(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net511),
    .X(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net783),
    .S(net323),
    .X(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[68] ),
    .Y(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1  (.A1(net400),
    .A2(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net266),
    .X(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y  (.A(net473),
    .B(net477),
    .Y(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[69] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[69] ),
    .A1(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net518),
    .X(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net746),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B  (.A(net494),
    .B(\m_blake2.m_hash256.h_flat[69] ),
    .X(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1  (.A1(net288),
    .A2(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net283),
    .C1(net354),
    .X(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[70] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[70] ),
    .A1(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net854),
    .S(net332),
    .X(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[70] ),
    .Y(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22ai_1 \m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2  (.A1(net266),
    .A2(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B2(net400),
    .Y(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[71] ),
    .X(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net281),
    .A2(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(net355),
    .X(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[71] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[71] ),
    .A1(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net670),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[72] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[72] ),
    .A1(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net757),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B  (.A(net486),
    .B(\m_blake2.m_hash256.h_flat[72] ),
    .Y(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1  (.A1(net400),
    .A2(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net266),
    .C1(net366),
    .X(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[73] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[73] ),
    .A1(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net501),
    .X(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net909),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[73] ),
    .X(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B  (.A(net277),
    .B(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__and2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[74] ),
    .X(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[74] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[74] ),
    .A1(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net689),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[75] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[75] ),
    .A1(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net528),
    .X(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net840),
    .S(net335),
    .X(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__nand2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[75] ),
    .Y(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[76] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[76] ),
    .A1(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net511),
    .X(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net915),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B  (.A(net489),
    .B(\m_blake2.m_hash256.h_flat[76] ),
    .X(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1  (.A1(net285),
    .A2(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net279),
    .C1(net350),
    .X(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[77] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[77] ),
    .A1(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net518),
    .X(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net724),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[77] ),
    .X(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2  (.A1(net283),
    .A2(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net288),
    .C1(net354),
    .X(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[78] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[78] ),
    .A1(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net781),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[78] ),
    .Y(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22ai_1 \m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2  (.A1(net266),
    .A2(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net400),
    .Y(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[79] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[79] ),
    .A1(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net862),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B  (.A(net495),
    .B(\m_blake2.m_hash256.h_flat[79] ),
    .Y(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2  (.A1(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ),
    .A2(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net400),
    .X(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[80] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[80] ),
    .A1(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net817),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[80] ),
    .Y(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B  (.A(net266),
    .B(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nand2_4 \m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y  (.A(net473),
    .B(net407),
    .Y(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[81] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[81] ),
    .A1(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net502),
    .X(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net710),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[81] ),
    .X(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N  (.A1_N(net277),
    .A2_N(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net400),
    .X(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[82] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[82] ),
    .A1(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net660),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[82] ),
    .X(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N  (.A1_N(net277),
    .A2_N(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(net400),
    .X(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[83] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[83] ),
    .A1(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net528),
    .X(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net790),
    .S(net334),
    .X(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[83] ),
    .X(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net281),
    .A2(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net287),
    .X(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[84] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[84] ),
    .A1(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net510),
    .X(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net789),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__nand2_2_B  (.A(net434),
    .B(\m_blake2.m_hash256.h_flat[84] ),
    .Y(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[85] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[85] ),
    .A1(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net755),
    .S(net324),
    .X(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[85] ),
    .X(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2  (.A1(net283),
    .A2(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .C1(net354),
    .Y(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[86] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[86] ),
    .A1(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net830),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B  (.A(net497),
    .B(\m_blake2.m_hash256.h_flat[86] ),
    .Y(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2  (.A1(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ),
    .A2(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ),
    .C1(net389),
    .X(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[87] ),
    .X(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net280),
    .A2(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .X(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[87] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[87] ),
    .A1(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net681),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B  (.A(net434),
    .B(\m_blake2.m_hash256.h_flat[88] ),
    .X(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net279),
    .A2(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ),
    .C1(net350),
    .X(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[88] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[88] ),
    .A1(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net1737),
    .S(net318),
    .X(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[89] ),
    .X(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net278),
    .A2(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_Y ),
    .C1(net346),
    .X(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[89] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[89] ),
    .A1(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net502),
    .X(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net884),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(net731),
    .S(net309),
    .X(\m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[8] ),
    .A1(\m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net502),
    .X(\hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__mux2_1_A0_A1_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C_X ),
    .B(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .Y(\m_blake2.m_hash256.h_flat[8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[90] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[90] ),
    .A1(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net793),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B  (.A(net483),
    .B(\m_blake2.m_hash256.h_flat[90] ),
    .X(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net277),
    .A2(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net289),
    .X(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[91] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[91] ),
    .A1(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net528),
    .X(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net743),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[91] ),
    .X(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net280),
    .A2(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net287),
    .X(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[92] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[92] ),
    .A1(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net510),
    .X(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net888),
    .S(net326),
    .X(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B  (.A(net490),
    .B(\m_blake2.m_hash256.h_flat[92] ),
    .Y(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2  (.A1(net266),
    .A2(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2 ),
    .X(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .B(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ),
    .Y(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[93] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[93] ),
    .A1(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net517),
    .X(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net896),
    .S(net325),
    .X(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B  (.A(net494),
    .B(\m_blake2.m_hash256.h_flat[93] ),
    .Y(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2  (.A1(net266),
    .A2(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ),
    .X(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B  (.A(net437),
    .B(\m_blake2.m_hash256.h_flat[94] ),
    .X(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(net286),
    .A2(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net280),
    .X(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[94] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[94] ),
    .A1(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net525),
    .X(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net706),
    .S(net331),
    .X(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B  (.A(net438),
    .B(\m_blake2.m_hash256.h_flat[95] ),
    .X(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net280),
    .A2(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net287),
    .X(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[95] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[95] ),
    .A1(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net526),
    .X(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net709),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B  (.A(net429),
    .B(\m_blake2.m_hash256.h_flat[96] ),
    .X(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net284),
    .A2(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(net346),
    .X(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[96] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[96] ),
    .A1(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net511),
    .X(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net857),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[97] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[97] ),
    .A1(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net505),
    .X(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net715),
    .S(net313),
    .X(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B  (.A(net484),
    .B(\m_blake2.m_hash256.h_flat[97] ),
    .X(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2  (.A1(net284),
    .A2(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__or2_2_B_X ),
    .B2(net277),
    .C1(net346),
    .X(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__and2_2_B  (.A(net428),
    .B(\m_blake2.m_hash256.h_flat[98] ),
    .X(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[98] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[98] ),
    .A1(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net750),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[99] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[99] ),
    .A1(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net527),
    .X(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A1(net695),
    .S(net333),
    .X(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B  (.A(net496),
    .B(\m_blake2.m_hash256.h_flat[99] ),
    .X(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2  (.A1(net287),
    .A2(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__and2_2_B_X ),
    .B2(net280),
    .C1(net359),
    .X(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.h_flat[9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ),
    .A1(net703),
    .S(net311),
    .X(\m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.h_flat[9] ),
    .A1(\m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net503),
    .X(\hash[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.last_block_q ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.last_block_q ),
    .B(net344),
    .Y(\m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[0] ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2 ),
    .B1_N(\m_blake2.m_hash256.g_b[0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2 ));
 sky130_fd_sc_hd__or3_2 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X  (.A(net106),
    .B(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B ),
    .C(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][0] ),
    .A2(net98),
    .B1(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1 ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][0] ),
    .A2(net110),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][0] ),
    .A2(net114),
    .B1(net138),
    .B2(\m_blake2.m_hash256.m_matrix[2][0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][0] ),
    .A2(net126),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][0] ),
    .A2(net86),
    .B1(net130),
    .B2(\m_blake2.m_hash256.m_matrix[8][0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][0] ),
    .A2(net146),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][0] ),
    .A2(net134),
    .B1(net118),
    .B2(\m_blake2.m_hash256.m_matrix[13][0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][0] ),
    .A2(net90),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][0] ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[10] ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .B(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[11] ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a31o_2_X  (.A1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .A3(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .X(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .A2(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[12] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__a311oi_4 \m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a311oi_2_Y  (.A1(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.a0[10]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .A3(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B ),
    .C1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[13] ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[14] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or3_2_B  (.A(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .C(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__o311a_1 \m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o311a_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A3(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[13]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .C1(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[15] ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .B(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__a31oi_4 \m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2  (.A1(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .A3(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .Y(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[16] ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ),
    .C(\m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .X(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__nor3_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__nor3_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ),
    .C(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[17] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2_Y ),
    .B1(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[17]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[18] ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_A_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .A2(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .B1(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_A ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .C(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .Y(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2_Y ),
    .B(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .Y(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[19] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3  (.A1(\m_blake2.m_hash256.m_g.a0[15]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a31oi_2_A2_Y ),
    .A2(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .A3(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a221o_2_C1_X ),
    .X(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a0[18]_sky130_fd_sc_hd__and2_2_X_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[1] ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__or3b_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .C_N(\m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__or3b_2_X_C_N ),
    .X(\m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3_X ),
    .X(\m_blake2.m_hash256.m_g.a0[20] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[21] ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_Y ),
    .B(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21bo_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B1_N(\m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21bo_2_X_B1_N ),
    .X(\m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[22] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3_X ),
    .A2(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .B1(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_Y ),
    .B(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.m_g.a0[20]_sky130_fd_sc_hd__xor2_2_X_A ),
    .X(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[21]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21bo_2_X_B1_N ),
    .A2(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_Y ),
    .B1(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[23] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A3 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[24] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .B(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[19]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__a31o_2_A3_X ),
    .A2(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .A3(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A3 ),
    .B1(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1 ),
    .X(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .A2(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A3 ),
    .B1(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_g.a0[23]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a31o_2_X_B1 ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[25] ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_A_N ),
    .B(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_A_N_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .B(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_A_N ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ),
    .B(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[26] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a31oi_2 \m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[24]_sky130_fd_sc_hd__and2_2_X_A ),
    .A3(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_A_N ),
    .Y(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[27] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ),
    .A2(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .B(\m_blake2.m_hash256.m_g.a0[26]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[28] ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X  (.A1_N(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A ),
    .A2_N(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X ),
    .B2(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2 ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__o32a_4 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net101),
    .B2(\m_blake2.m_hash256.m_matrix[0][27] ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][27] ),
    .A2(net91),
    .B1(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net107),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][27] ),
    .A2(net147),
    .B1(net151),
    .B2(\m_blake2.m_hash256.m_matrix[11][27] ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][27] ),
    .A2(net126),
    .B1(net139),
    .B2(\m_blake2.m_hash256.m_matrix[2][27] ),
    .C1(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][27] ),
    .A2(net87),
    .B1(net119),
    .B2(\m_blake2.m_hash256.m_matrix[13][27] ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][27] ),
    .A2(net111),
    .B1(net114),
    .B2(\m_blake2.m_hash256.m_matrix[5][27] ),
    .C1(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][27] ),
    .A2(net95),
    .B1(net123),
    .B2(\m_blake2.m_hash256.m_matrix[15][27] ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][27] ),
    .A2(net134),
    .B1(net143),
    .B2(\m_blake2.m_hash256.m_matrix[1][27] ),
    .C1(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][27] ),
    .A2(net131),
    .B1(net99),
    .B2(\m_blake2.m_hash256.m_matrix[6][27] ),
    .X(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .A2(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[29] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__nor3_2_Y  (.A(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_X ),
    .C(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[2] ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21ba_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1_N(\m_blake2.m_hash256.m_g.a0[1]_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__or3b_2_X_C_N ),
    .X(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .B(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_A_N_sky130_fd_sc_hd__o21ba_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__or3b_2_X_A ),
    .A2(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1_N(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_A_N ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__or3b_2_X  (.A(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__or3b_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_X ),
    .C_N(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[30] ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__o21ba_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1_N(\m_blake2.m_hash256.m_g.a0[29]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[31] ));
 sky130_fd_sc_hd__o21bai_1 \m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21bai_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1_N(\m_blake2.m_hash256.m_g.a0[30]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__or2_2_X_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_Y ),
    .B(\m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[31]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[3] ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .B(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_X ),
    .X(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_X ),
    .B(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .X(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[4] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .A2(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[3]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .X(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[5] ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_X ),
    .X(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_B1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[6] ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .B(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_A_N_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .A2(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X  (.A(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_A ),
    .B(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_X ),
    .C_N(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_C_N ),
    .X(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[4]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ),
    .C1(\m_blake2.m_hash256.m_g.a0[5]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[7] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X  (.A1(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B ),
    .A3(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_A_N ),
    .X(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.a0[8] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .B(\m_blake2.m_hash256.m_g.a0[7]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[9] ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y  (.A1(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.a0[8]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ),
    .X(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.a0[9]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__a21o_2 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[0] ),
    .A2(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__a31o_2 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A3(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X ));
 sky130_fd_sc_hd__a21o_2 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.m_g.a0[0] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[0] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[0] ),
    .B(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__a21oi_4 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[10] ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__and2b_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a311o_1 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1  (.A1(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .A3(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21boi_2_B1_N_Y ),
    .C1(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__and3b_2_A_N_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__and3b_2_A_N_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1_A2 ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.m_g.a0[10] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[10] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[10] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.m_g.a0[11] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[11] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[11] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[12] ),
    .B(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.m_g.a0[12] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[12] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[12] ),
    .B(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__o21bai_2 \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1_A2 ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.m_g.a0[13] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[13] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[13] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[13] ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__o31a_2 \m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o31a_2_B1_A2 ),
    .A3(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2 ));
 sky130_fd_sc_hd__a21oi_4 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[14] ),
    .A2(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.m_g.a0[14] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[14] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[14] ),
    .B(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2 ),
    .B1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2 ),
    .X(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21a_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_4 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[15] ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.m_g.a0[15] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[15] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[15] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__o311a_1 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1  (.A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .A3(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C1(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nor4_2 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D  (.A(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .D(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a311o_2_C1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A1 ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y_sky130_fd_sc_hd__nand3_2_C  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__and3b_2_A_N_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A2 ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[16] ),
    .A2(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.m_g.a0[16] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[16] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[16] ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A ),
    .A2(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_A1 ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A1 ),
    .A2(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A2 ),
    .A3(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_A1 ));
 sky130_fd_sc_hd__or4bb_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ),
    .C_N(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ),
    .D_N(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A1 ),
    .A2(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a31o_2_B1_A2 ),
    .A3(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a21bo_2 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X  (.A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1 ),
    .A2(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor4_2_D_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o311a_2_C1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1 ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.m_g.a0[17] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[17] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[17] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[18] ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_C ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.m_g.a0[18] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[18] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[18] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__nand3_2 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B1(\m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand3_2_B  (.A(\m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_A1 ),
    .A2(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__or3_2 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__o21bai_4 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__o21bai_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_A1 ),
    .A2(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.m_g.a0[19] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[19] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.m_g.a0[1] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[1] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[1] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o21bai_1 \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_X ),
    .B1_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[20] ),
    .A2(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A2 ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.m_g.a0[20] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[20] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[20] ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[21] ),
    .A2(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A2 ),
    .Y(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.m_g.a0[21] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[21] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[21] ),
    .B(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.m_g.a0[22] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[22] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[22] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[22] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A2 ),
    .B1(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B2(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X ));
 sky130_fd_sc_hd__a31oi_2 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21ba_2_A2_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ),
    .A3(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.m_g.a0[23] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[23] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[23] ),
    .B(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[23] ),
    .B(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.m_g.a0[24] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[24] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[24] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[24] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a21oi_4 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X_sky130_fd_sc_hd__a31o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or4bb_2_A_X_sky130_fd_sc_hd__a31o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__a31oi_2_B1_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.m_g.a0[25] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[25] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[25] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.m_g.a0[26] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[26] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[26] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.m_g.a0[27] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[27] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[27] ),
    .B(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[27] ),
    .B(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[28] ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.m_g.a0[28] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[28] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[28] ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__o211ai_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C1(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y ));
 sky130_fd_sc_hd__o311a_4 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A3(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y ),
    .C1(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_B1 ),
    .X(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_B1 ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[29] ),
    .A2(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.m_g.a0[29] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[29] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[29] ),
    .B(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__o21bai_1 \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y ));
 sky130_fd_sc_hd__o311a_2 \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A3(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_B1 ),
    .C1(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_X ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_X ),
    .C_N(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3b_2_C_N_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.m_g.a0[2] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[2] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[2] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21bai_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[30] ),
    .A2(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_50_clk),
    .D(\m_blake2.m_hash256.m_g.a0[30] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[30] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[30] ),
    .B(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_50_clk),
    .D(\m_blake2.m_hash256.m_g.a0[31] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[31] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.m_g.a0[3] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[3] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[3] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__and3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ba_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ba_2_A1_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__and3_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .C(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[4] ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_63_clk),
    .D(\m_blake2.m_hash256.m_g.a0[4] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[4] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[4] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ba_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_A2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ba_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ba_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.a_q[5] ),
    .X(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .A3(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_A2 ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_A2 ),
    .Y(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[5] ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_C ),
    .X(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_B ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_63_clk),
    .D(\m_blake2.m_hash256.m_g.a0[5] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[5] ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[6] ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_63_clk),
    .D(\m_blake2.m_hash256.m_g.a0[6] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[6] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[6] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nor3b_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_A ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_X ),
    .C_N(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y ));
 sky130_fd_sc_hd__a21boi_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a31o_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y ),
    .A3(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a31o_2_A2_X ));
 sky130_fd_sc_hd__and3_2 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y ),
    .C(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_A ),
    .A2(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__and3_2_A_X ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .B2(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C1(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and3b_2_B_X_sky130_fd_sc_hd__a31o_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_B1_N_X_sky130_fd_sc_hd__a221o_2_B1_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_63_clk),
    .D(\m_blake2.m_hash256.m_g.a0[7] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[7] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[7] ),
    .Y(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__and3_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__or3_2 \m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__and3_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.m_g.a0[8] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[8] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[8] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[8] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.m_g.a0[9] ),
    .Q(\m_blake2.m_hash256.m_g.a_q[9] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[9] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__a21boi_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21boi_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21boi_2_B1_N_Y ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[9] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__and3b_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__and3b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__and3b_2_A_N_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a31o_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__o31a_2 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__and3_2_B_X ),
    .A3(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_b[0] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[0] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[0] ),
    .B(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand2_4 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.g_b[10] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[10] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[10] ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_1  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1 ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B1(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[11] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[11] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[11] ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2  (.A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1 ),
    .A2(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .A3(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B2(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1 ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1 ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o41a_2_B1_A3 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__o41a_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o41a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X ),
    .A3(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o41a_2_B1_A3 ),
    .A4(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_C ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_C ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X ),
    .C_N(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__or3b_2_B_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[31]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_b[12] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[12] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[12] ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A3(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__o21ai_4 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2  (.A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__or4bb_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__or4bb_2_C_N  (.A(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .C_N(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X ),
    .D_N(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__or4bb_2_C_N_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .A2(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .C(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__o21bai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .D(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__o2111a_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2  (.A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__or4bb_2_C_N_X ),
    .C1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .D1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_b[13] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[13] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[13] ),
    .Y(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand3_2 \m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.b_q[14] ),
    .X(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_b[14] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[14] ));
 sky130_fd_sc_hd__nand3_2 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[14] ),
    .B(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .C(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .B1(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .C(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y_C_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .A2(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .C1(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y_C ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.b_q[15] ),
    .X(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[15] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[15] ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[15] ),
    .B(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .C(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_63_clk),
    .D(\m_blake2.m_hash256.g_b[16] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[16] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16] ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C  (.A(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .D(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .D(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or4_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .D(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_A2 ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_B ),
    .C(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__o21bai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.b_q[17] ),
    .X(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.g_b[17] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[17] ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[17] ),
    .B(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .X(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X_B1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_C ),
    .X(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .C(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__a21o_2_X_B1 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_C ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.g_b[18] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[18] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[18] ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a2111o_2_A2  (.A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .C1(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .D1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a2111o_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__or4_2_C_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__a31o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .A3(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.b_q[19] ),
    .X(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.g_b[19] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[19] ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[19] ),
    .B(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .C(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.g_b[1] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[1] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[1] ),
    .B(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.g_b[20] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[20] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[20] ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_B1 ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2 ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_B1_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_B1 ));
 sky130_fd_sc_hd__o21a_2 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_B ),
    .B1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__and2_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ),
    .B1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__and2_2_B_X ),
    .C(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[21] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[21] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[21] ),
    .B(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[22] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[22] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[22] ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__o21bai_2 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[23] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[23] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[23] ),
    .B(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2  (.A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A3(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B2(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__o211a_2 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o2111a_2_A2_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_A2 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X ),
    .C1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a2111o_2_A2_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[24] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[24] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[24] ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .C(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A1 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A1 ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A1 ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.g_b[25] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[25] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[25] ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__a21o_2 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_A1 ),
    .A2(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2  (.A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_A1 ),
    .A2(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_A1_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_A1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_A1 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o32a_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .A3(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3 ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1_sky130_fd_sc_hd__a21o_2_A2  (.A1(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1 ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B_A ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_B1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_A3 ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_b[26] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[26] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[26] ),
    .B(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_b[27] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[27] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[27] ),
    .B(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[28] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[28] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[28] ),
    .B(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_A ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .X(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .B1(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_50_clk),
    .D(\m_blake2.m_hash256.g_b[29] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[29] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[29] ),
    .B(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[17]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_b[2] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[2] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[2] ),
    .B(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_B1 ),
    .B(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B2 ),
    .B(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_50_clk),
    .D(\m_blake2.m_hash256.g_b[30] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[30] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[30] ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a32o_2 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2  (.A1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1 ),
    .A2(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .A3(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3 ),
    .B1(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B2(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1 ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1 ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3 ));
 sky130_fd_sc_hd__o21bai_4 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2_sky130_fd_sc_hd__o21bai_2_Y  (.A1(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o211a_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or3_2_B_X ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__o32a_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X ),
    .B(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X  (.A(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2 ),
    .A3(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_2 \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[31] ),
    .X(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.g_b[31] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[31] ));
 sky130_fd_sc_hd__nand3b_4 \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[31] ),
    .B(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y ),
    .C(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_b[3] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[3] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[3] ),
    .B(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a21oi_4 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_49_clk),
    .D(\m_blake2.m_hash256.g_b[4] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[4] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[4] ),
    .B(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__and2b_2 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N ),
    .B(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_B ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2  (.A1(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_b[5] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[5] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[5] ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__o31ai_4 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__o31ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .A3(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_A2 ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21ba_2_A2_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[25]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2_B1 ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.g_b[6] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[6] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[6] ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__o31ai_4 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_A2 ),
    .A3(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_B1 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_A2 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_A2 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .B1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_B1 ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_b[7] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[7] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[7] ),
    .B(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_64_clk),
    .D(\m_blake2.m_hash256.g_b[8] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[8] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[8] ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__o21bai_2 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__o41a_2_B1_A3 ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__o31ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__o21bai_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_X ),
    .C(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.g_b[9] ),
    .Q(\m_blake2.m_hash256.m_g.b_q[9] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[9] ),
    .B(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.g_c[0] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[0] ));
 sky130_fd_sc_hd__nand2_4 \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[0] ),
    .B(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[0] ),
    .B(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a41o_2 \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2  (.A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A4(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X ));
 sky130_fd_sc_hd__a21bo_4 \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B1_N(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X ),
    .B(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.g_c[10] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[10] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[10] ),
    .B(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B ),
    .B1(\m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[10] ),
    .B(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[11] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_B1 ),
    .Y(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_c[11] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[11] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[11] ),
    .B(\m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__o22ai_1 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o22ai_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[11] ),
    .B(\m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__or4_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__or3_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .D(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_A4 ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__a21o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[12] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B2(\m_blake2.m_hash256.m_g.c_q[13] ),
    .X(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.g_c[12] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[12] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[12] ),
    .B(\m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B1(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__nand3_2 \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .C(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[12] ),
    .B(\m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.g_c[13] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[13] ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[13] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_C_sky130_fd_sc_hd__nand3_2_Y_C ),
    .B1(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_A4 ),
    .X(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_B ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[13] ),
    .B(\m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_c[14] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[14] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[14] ),
    .B(\m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[14] ),
    .B(\m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[15] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__o211a_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__o41a_1 \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[12]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[11]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .A3(\m_blake2.m_hash256.m_g.c_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A4(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_A4 ),
    .B1(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_X ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_X_sky130_fd_sc_hd__a31o_2_A3  (.A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_B ),
    .A3(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.g_c[15] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[15] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__o211a_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[15] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X ),
    .C1(\m_blake2.m_hash256.m_g.c_q[14] ),
    .X(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__o211a_2_A1_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[15] ),
    .B(\m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[14]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_A4 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.g_c[16] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[16] ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[16] ),
    .B(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[16] ),
    .B(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_B ),
    .A3(\m_blake2.m_hash256.m_g.c_q[15]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__o41a_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_B ),
    .C(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A_Y ),
    .D(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__nand2b_2_Y  (.A_N(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.g_c[17] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[17] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[17] ),
    .B(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[17] ),
    .B(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.g_c[18] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[18] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[18] ),
    .B(\m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[18] ),
    .B(\m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a311o_1 \m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a311o_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .A3(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C1(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand3_2_Y_B ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[19] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B2 ),
    .C1(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__o211a_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1 ),
    .Y(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.m_g.c_q[18]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B2_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B2 ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__o31a_2 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o31a_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or4_2_A_B ),
    .A3(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__inv_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.g_c[19] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[19] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__o211a_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[19] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .C1(\m_blake2.m_hash256.m_g.c_q[18] ),
    .X(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__o211a_2_A1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[19] ),
    .B(\m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.g_c[1] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[1] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[1] ),
    .B(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B2 ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[1] ),
    .B(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[1]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[20] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B2(\m_blake2.m_hash256.m_g.c_q[21] ),
    .X(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_63_clk),
    .D(\m_blake2.m_hash256.g_c[20] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[20] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[20] ),
    .B(\m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[20] ),
    .B(\m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.g_c[21] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[21] ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[21] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__o21ai_2_A1_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ),
    .A2(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[21] ),
    .B(\m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[20]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_c[22] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[22] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[22] ),
    .B(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .B1(\m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[22] ),
    .B(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_c[23] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[23] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[23] ),
    .B(\m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[23] ),
    .B(\m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2  (.A1(\m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .C1(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[23] ),
    .B(\m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[23]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.g_c[24] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[24] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[24] ),
    .B(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[24] ),
    .B(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_B ),
    .A2(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_C ),
    .B1(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .C(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.g_c[25] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[25] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[25] ),
    .B(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[25] ),
    .B(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2  (.A1(\m_blake2.m_hash256.m_g.c_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__o21a_2 \m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A2(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.g_c[26] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[26] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[26] ),
    .B(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[26] ),
    .B(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_c[27] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[27] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[27] ),
    .B(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[27] ),
    .B(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2  (.A1(\m_blake2.m_hash256.m_g.c_q[26]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.m_g.c_q[25]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C1(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A2(\m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__o221a_2_A2_X ),
    .B1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_63_clk),
    .D(\m_blake2.m_hash256.g_c[28] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[28] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[28] ),
    .B(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[28] ),
    .B(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_c[29] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[29] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[29] ),
    .B(\m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[29] ),
    .B(\m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[2] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_B1 ),
    .Y(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and2b_2_X  (.A_N(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B2 ),
    .X(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__a21oi_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.g_c[2] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[2] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[2] ),
    .B(\m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_c[30] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[30] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[30] ),
    .B(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[30] ),
    .B(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.g_c[31] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[31] ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[31] ),
    .B(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_B ),
    .B1(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__nand3_2 \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C  (.A(\m_blake2.m_hash256.m_g.c_q[30]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_B ),
    .C(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y ));
 sky130_fd_sc_hd__a311o_1 \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_B_sky130_fd_sc_hd__a311o_2_X  (.A1(\m_blake2.m_hash256.m_g.c_q[28]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a31o_2_X_A2 ),
    .A3(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[29]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .C1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A ),
    .X(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_B ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .Y(\m_blake2.m_hash256.m_g.c_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a221oi_4 \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[3] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B2 ),
    .C1(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__o211a_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.g_c[3] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[3] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__o211a_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[3] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .C1(\m_blake2.m_hash256.m_g.c_q[2] ),
    .X(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__o211a_2_A1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[3] ),
    .B(\m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.g_c[4] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[4] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[4] ),
    .B(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[4] ),
    .B(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.g_c[5] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[5] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[5] ),
    .B(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[5] ),
    .B(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__o21a_2 \m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N ),
    .B1(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_c[6] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[6] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[6] ),
    .B(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_A_B ),
    .X(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[6] ),
    .B(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.g_c[7] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[7] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[7] ),
    .B(\m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1  (.A1(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_A2 ),
    .B1(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_B1 ),
    .C1(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_X ));
 sky130_fd_sc_hd__o21bai_2 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__o21bai_2_A1  (.A1(\m_blake2.m_hash256.m_g.c_q[7] ),
    .A2(\m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B1_N(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__o21bai_2_A1_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[7] ),
    .B(\m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand3b_1 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__or2_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.c_q[5]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_B1 ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .C(\m_blake2.m_hash256.m_g.c_q[4]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.g_c[8] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[8] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[8] ),
    .B(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .Y(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[8] ),
    .B(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__o21bai_2_A1_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_X ),
    .B1(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.g_c[9] ),
    .Q(\m_blake2.m_hash256.m_g.c_q[9] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[9] ),
    .B(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.c_q[9] ),
    .B(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.m_g.c_q[8]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.c_q[9]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_d[0] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[0] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[0] ),
    .B(\m_blake2.m_hash256.m_g.a_q[0] ),
    .X(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_d[10] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[10] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[10] ),
    .B(\m_blake2.m_hash256.m_g.d_q[10] ),
    .X(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.g_d[11] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[11] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[11] ),
    .B(\m_blake2.m_hash256.m_g.d_q[11] ),
    .X(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.g_d[12] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[12] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[12] ),
    .B(\m_blake2.m_hash256.m_g.d_q[12] ),
    .X(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .X(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_d[13] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[13] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[13] ),
    .B(\m_blake2.m_hash256.m_g.d_q[13] ),
    .X(\m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.g_d[14] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[14] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[14] ),
    .B(\m_blake2.m_hash256.m_g.d_q[14] ),
    .X(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_50_clk),
    .D(\m_blake2.m_hash256.g_d[15] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[15] ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[15] ),
    .B(\m_blake2.m_hash256.m_g.d_q[15] ),
    .Y(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.g_d[16] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[16] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[16] ),
    .B(\m_blake2.m_hash256.m_g.a_q[16] ),
    .X(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_d[17] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[17] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[17] ),
    .B(\m_blake2.m_hash256.m_g.a_q[17] ),
    .X(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_d[18] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[18] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[18] ),
    .B(\m_blake2.m_hash256.m_g.a_q[18] ),
    .X(\m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_d[19] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[19] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[19] ),
    .B(\m_blake2.m_hash256.m_g.a_q[19] ),
    .X(\m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_d[1] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[1] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[1] ),
    .B(\m_blake2.m_hash256.m_g.a_q[1] ),
    .X(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_d[20] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[20] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[20] ),
    .B(\m_blake2.m_hash256.m_g.a_q[20] ),
    .X(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_d[21] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[21] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[21] ),
    .B(\m_blake2.m_hash256.m_g.a_q[21] ),
    .X(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_d[22] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[22] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[22] ),
    .B(\m_blake2.m_hash256.m_g.a_q[22] ),
    .X(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_50_clk),
    .D(\m_blake2.m_hash256.g_d[23] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[23] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[23] ),
    .B(\m_blake2.m_hash256.m_g.a_q[23] ),
    .X(\m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_d[24] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[24] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[24] ),
    .B(\m_blake2.m_hash256.m_g.a_q[24] ),
    .X(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.g_d[25] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[25] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[25] ),
    .B(\m_blake2.m_hash256.m_g.a_q[25] ),
    .X(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.g_d[26] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[26] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[26] ),
    .B(\m_blake2.m_hash256.m_g.a_q[26] ),
    .X(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_d[27] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[27] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[27] ),
    .B(\m_blake2.m_hash256.m_g.a_q[27] ),
    .X(\m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.g_d[28] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[28] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[28] ),
    .B(\m_blake2.m_hash256.m_g.a_q[28] ),
    .X(\m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_d[29] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[29] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[29] ),
    .B(\m_blake2.m_hash256.m_g.a_q[29] ),
    .X(\m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.g_d[2] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[2] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[2] ),
    .B(\m_blake2.m_hash256.m_g.a_q[2] ),
    .X(\m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_d[30] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[30] ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[30] ),
    .B(\m_blake2.m_hash256.m_g.a_q[30] ),
    .X(\m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.g_d[31] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[31] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[31] ),
    .B(\m_blake2.m_hash256.m_g.a_q[31] ),
    .X(\m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.g_d[3] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[3] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[3] ),
    .B(\m_blake2.m_hash256.m_g.a_q[3] ),
    .X(\m_blake2.m_hash256.m_g.d_q[3]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.g_d[4] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[4] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[4] ),
    .B(\m_blake2.m_hash256.m_g.a_q[4] ),
    .X(\m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.g_d[5] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[5] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[5] ),
    .B(\m_blake2.m_hash256.m_g.a_q[5] ),
    .X(\m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.g_d[6] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[6] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[6] ),
    .B(\m_blake2.m_hash256.m_g.d_q[6] ),
    .X(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.g_d[7] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[7] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[7] ),
    .B(\m_blake2.m_hash256.m_g.d_q[7] ),
    .X(\m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .X(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.g_d[8] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[8] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[8] ),
    .B(\m_blake2.m_hash256.m_g.d_q[8] ),
    .X(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.g_d[9] ),
    .Q(\m_blake2.m_hash256.m_g.d_q[9] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[9] ),
    .B(\m_blake2.m_hash256.m_g.d_q[9] ),
    .X(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.g_y[0] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.g_y[10] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10] ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10] ),
    .B(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.g_y[11] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11] ),
    .B(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o21a_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[11]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__xnor2_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11] ),
    .B(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12] ),
    .B(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[12]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.g_y[12] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12] ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.g_y[13] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[13] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[13] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.g_y[14] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15] ),
    .B(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.g_y[15] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15] ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15] ),
    .B(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16] ),
    .B(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.g_y[16] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.g_y[17] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.g_y[18] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18] ),
    .B(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N  (.A1(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ),
    .A2(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .B1_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[19] ),
    .X(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__nand3_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[19] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .C(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__and3_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.g_y[19] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19] ));
 sky130_fd_sc_hd__nand3b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19] ),
    .B(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ),
    .C(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__a21bo_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[19] ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.g_y[1] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.g_y[20] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21] ),
    .B(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.g_y[21] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21] ),
    .B(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.g_y[22] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22] ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21o_2_A1_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22] ),
    .B(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.g_y[23] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23] ),
    .B(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23] ),
    .B(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.g_y[24] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24] ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2_B1 ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a21boi_4 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2  (.A1(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .B1_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nand3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_C ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__o221a_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2  (.A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_A1_X ),
    .A2(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2_B1 ),
    .B2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y ),
    .C1(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o221a_2_B2_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .A2(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__xnor2_4 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24] ),
    .B(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.g_y[25] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25] ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.g_y[26] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26] ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26] ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.g_y[27] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27] ),
    .B(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27] ),
    .B(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28] ),
    .B(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_B_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_A_N_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.g_y[28] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29] ),
    .B(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_4 \m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.g_y[29] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29] ),
    .B(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2] ),
    .B(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.g_y[2] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[2] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.g_y[30] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.g_y[31] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[31] ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[31]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.m_g.a_q[31] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[31] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[31]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3] ),
    .B(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.g_y[3] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3] ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.g_y[4] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4] ),
    .B(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.g_y[5] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5] ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_A ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6] ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.g_y[6] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6] ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6] ),
    .B(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .A2(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .B1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ),
    .B(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .C(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.g_y[7] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_X  (.A(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B ),
    .B(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.a_q[7]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__or3_2_A_X ),
    .C(\m_blake2.m_hash256.m_g.a_q[8]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.g_y[8] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8] ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8] ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8] ),
    .B(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.g_y[9] ),
    .Q(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9] ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9] ),
    .B(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9] ),
    .B(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net769),
    .A1(\m_blake2.m_hash256.m_matrix[0][8] ),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][0] ),
    .B(net103),
    .X(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2 ),
    .C(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1088),
    .A1(\m_blake2.m_hash256.m_matrix[0][18] ),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(net1319),
    .Q(\m_blake2.m_hash256.m_matrix[0][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1318),
    .A1(\m_blake2.m_hash256.m_matrix[0][19] ),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[0][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1121),
    .A1(\m_blake2.m_hash256.m_matrix[0][20] ),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[0][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][13] ),
    .A1(net1529),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[0][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1487),
    .A1(net1310),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[0][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(net1545),
    .Q(\m_blake2.m_hash256.m_matrix[0][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1544),
    .A1(\m_blake2.m_hash256.m_matrix[0][23] ),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[0][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1639),
    .A1(\m_blake2.m_hash256.m_matrix[0][24] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1143),
    .A1(net986),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[0][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][18] ),
    .A1(net1118),
    .S(net602),
    .X(\m_blake2.m_hash256.m_matrix[0][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1437),
    .A1(\m_blake2.m_hash256.m_matrix[0][27] ),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[0][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1094),
    .A1(\m_blake2.m_hash256.m_matrix[0][9] ),
    .S(net556),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2  (.A1(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1 ),
    .A2(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2 ),
    .A3(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3 ),
    .B1(net100),
    .B2(\m_blake2.m_hash256.m_matrix[0][1] ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][1] ),
    .A2(net110),
    .B1(net130),
    .B2(\m_blake2.m_hash256.m_matrix[8][1] ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][1] ),
    .A2(net90),
    .B1(net138),
    .B2(\m_blake2.m_hash256.m_matrix[2][1] ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][1] ),
    .A2(net86),
    .B1(net134),
    .B2(\m_blake2.m_hash256.m_matrix[3][1] ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][1] ),
    .A2(net118),
    .B1(net106),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][1] ),
    .A2(net146),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][1] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][1] ),
    .A2(net98),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][1] ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][1] ),
    .A2(net142),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][1] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][1] ),
    .A2(net126),
    .B1(net114),
    .B2(\m_blake2.m_hash256.m_matrix[5][1] ),
    .X(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X ),
    .B(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.m_g.a0[2]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__or3b_2_X_A ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X ),
    .B(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][20] ),
    .A1(\m_blake2.m_hash256.m_matrix[0][28] ),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[0][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(net1530),
    .Q(\m_blake2.m_hash256.m_matrix[0][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1529),
    .A1(\m_blake2.m_hash256.m_matrix[0][29] ),
    .S(net550),
    .X(\m_blake2.m_hash256.m_matrix[0][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1310),
    .A1(\m_blake2.m_hash256.m_matrix[0][30] ),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[0][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1868),
    .A1(\m_blake2.m_hash256.m_matrix[0][31] ),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[0][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][24] ),
    .A1(net1636),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[0][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net986),
    .A1(\m_blake2.m_hash256.m_matrix[1][1] ),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[0][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(net1119),
    .Q(\m_blake2.m_hash256.m_matrix[0][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1118),
    .A1(\m_blake2.m_hash256.m_matrix[1][2] ),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[0][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][27] ),
    .A1(net1899),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[0][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][28] ),
    .A1(\m_blake2.m_hash256.m_matrix[1][4] ),
    .S(net558),
    .X(\m_blake2.m_hash256.m_matrix[0][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1797),
    .A1(\m_blake2.m_hash256.m_matrix[1][5] ),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[0][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(net947),
    .Q(\m_blake2.m_hash256.m_matrix[0][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net946),
    .A1(\m_blake2.m_hash256.m_matrix[0][10] ),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2  (.A1(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1 ),
    .A2(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2 ),
    .A3(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3 ),
    .B1(net102),
    .B2(\m_blake2.m_hash256.m_matrix[0][2] ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][2] ),
    .A2(net110),
    .B1(net130),
    .B2(\m_blake2.m_hash256.m_matrix[8][2] ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][2] ),
    .A2(net115),
    .B1(net146),
    .B2(\m_blake2.m_hash256.m_matrix[10][2] ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][2] ),
    .A2(net87),
    .B1(net135),
    .B2(\m_blake2.m_hash256.m_matrix[3][2] ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][2] ),
    .A2(net139),
    .B1(net107),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][2] ),
    .A2(net98),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][2] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][2] ),
    .A2(net91),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][2] ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][2] ),
    .A2(net143),
    .B1(net95),
    .B2(\m_blake2.m_hash256.m_matrix[12][2] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][2] ),
    .A2(net127),
    .B1(net119),
    .B2(\m_blake2.m_hash256.m_matrix[13][2] ),
    .X(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X ),
    .Y(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A1_N ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X ),
    .B(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a2bb2o_2_B2_A2_N ),
    .Y(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][30] ),
    .A1(net1676),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[0][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][31] ),
    .A1(net1532),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[0][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(net871),
    .Q(\m_blake2.m_hash256.m_matrix[0][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net870),
    .A1(\m_blake2.m_hash256.m_matrix[0][11] ),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1  (.A1(\m_blake2.m_hash256.m_matrix[0][3] ),
    .A2(net102),
    .B1(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2 ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][3] ),
    .A2(net127),
    .B1(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net107),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][3] ),
    .A2(net134),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][3] ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][3] ),
    .A2(net86),
    .B1(net131),
    .B2(\m_blake2.m_hash256.m_matrix[8][3] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][3] ),
    .A2(net147),
    .B1(net123),
    .B2(\m_blake2.m_hash256.m_matrix[15][3] ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][3] ),
    .A2(net91),
    .B1(net99),
    .B2(\m_blake2.m_hash256.m_matrix[6][3] ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][3] ),
    .A2(net139),
    .B1(net151),
    .B2(\m_blake2.m_hash256.m_matrix[11][3] ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][3] ),
    .A2(net111),
    .B1(net115),
    .B2(\m_blake2.m_hash256.m_matrix[5][3] ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][3] ),
    .A2(net143),
    .B1(net118),
    .B2(\m_blake2.m_hash256.m_matrix[13][3] ),
    .X(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X ),
    .B(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_A2 ),
    .X(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.m_matrix[0][4] ),
    .A1(net1121),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22ai_4 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1  (.A1(\m_blake2.m_hash256.m_matrix[0][4] ),
    .A2(net100),
    .B1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2 ),
    .Y(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][4] ),
    .A2(net108),
    .B1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][4] ),
    .A2(net128),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][4] ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][4] ),
    .A2(net88),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][4] ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][4] ),
    .A2(net124),
    .B1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net104),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][4] ),
    .A2(net132),
    .B1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][4] ),
    .A2(net84),
    .B1(net96),
    .B2(\m_blake2.m_hash256.m_matrix[6][4] ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][4] ),
    .A2(net140),
    .B1(net116),
    .B2(\m_blake2.m_hash256.m_matrix[13][4] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][4] ),
    .A2(net112),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][4] ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][4] ),
    .A2(net136),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][4] ),
    .X(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__or3b_2_X_A ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X ),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.m_matrix[0][5] ),
    .A1(\m_blake2.m_hash256.m_matrix[0][13] ),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22ai_4 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1  (.A1(\m_blake2.m_hash256.m_matrix[0][5] ),
    .A2(net100),
    .B1(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2 ),
    .Y(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][5] ),
    .A2(net136),
    .B1(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net104),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][5] ),
    .A2(net112),
    .B1(net140),
    .B2(\m_blake2.m_hash256.m_matrix[1][5] ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][5] ),
    .A2(net108),
    .B1(net132),
    .B2(\m_blake2.m_hash256.m_matrix[3][5] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][5] ),
    .A2(net128),
    .B1(net96),
    .B2(\m_blake2.m_hash256.m_matrix[6][5] ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][5] ),
    .A2(net144),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][5] ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][5] ),
    .A2(net88),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][5] ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][5] ),
    .A2(net124),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][5] ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][5] ),
    .A2(net84),
    .B1(net116),
    .B2(\m_blake2.m_hash256.m_matrix[13][5] ),
    .X(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[6]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2b_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(net798),
    .Q(\m_blake2.m_hash256.m_matrix[0][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net797),
    .A1(\m_blake2.m_hash256.m_matrix[0][14] ),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1  (.A1(\m_blake2.m_hash256.m_matrix[0][6] ),
    .A2(net101),
    .B1(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2 ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][6] ),
    .A2(net145),
    .B1(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net105),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][6] ),
    .A2(net128),
    .B1(net93),
    .B2(\m_blake2.m_hash256.m_matrix[12][6] ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][6] ),
    .A2(net108),
    .B1(net121),
    .B2(\m_blake2.m_hash256.m_matrix[15][6] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][6] ),
    .A2(net117),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][6] ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][6] ),
    .A2(net132),
    .B1(net141),
    .B2(\m_blake2.m_hash256.m_matrix[1][6] ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][6] ),
    .A2(net137),
    .B1(net96),
    .B2(\m_blake2.m_hash256.m_matrix[6][6] ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][6] ),
    .A2(net84),
    .B1(net113),
    .B2(\m_blake2.m_hash256.m_matrix[5][6] ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][6] ),
    .A2(net125),
    .B1(net89),
    .B2(\m_blake2.m_hash256.m_matrix[14][6] ),
    .X(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X ),
    .B(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.m_matrix[0][7] ),
    .A1(net1544),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22ai_4 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1  (.A1(\m_blake2.m_hash256.m_matrix[0][7] ),
    .A2(net101),
    .B1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2 ),
    .Y(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][7] ),
    .A2(net89),
    .B1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][7] ),
    .A2(net141),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][7] ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][7] ),
    .A2(net133),
    .B1(net145),
    .B2(\m_blake2.m_hash256.m_matrix[10][7] ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][7] ),
    .A2(net137),
    .B1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net105),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][7] ),
    .A2(net125),
    .B1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][7] ),
    .A2(net85),
    .B1(net113),
    .B2(\m_blake2.m_hash256.m_matrix[5][7] ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][7] ),
    .A2(net129),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][7] ),
    .C1(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][7] ),
    .A2(net117),
    .B1(net93),
    .B2(\m_blake2.m_hash256.m_matrix[12][7] ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][7] ),
    .A2(net109),
    .B1(net97),
    .B2(\m_blake2.m_hash256.m_matrix[6][7] ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N  (.A_N(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .X(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y ),
    .B(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .Y(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][8] ),
    .A1(net1639),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[0][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[0][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[0][9] ),
    .A1(net1143),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(net1803),
    .Q(\m_blake2.m_hash256.m_matrix[10][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1802),
    .A1(\m_blake2.m_hash256.m_matrix[10][8] ),
    .S(net594),
    .X(\m_blake2.m_hash256.m_matrix[10][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(net1292),
    .Q(\m_blake2.m_hash256.m_matrix[10][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1291),
    .A1(\m_blake2.m_hash256.m_matrix[10][18] ),
    .S(net606),
    .X(\m_blake2.m_hash256.m_matrix[10][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1265),
    .A1(\m_blake2.m_hash256.m_matrix[10][19] ),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[10][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1091),
    .A1(\m_blake2.m_hash256.m_matrix[10][20] ),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[10][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1660),
    .A1(net1597),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[10][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1531),
    .A1(net1379),
    .S(net567),
    .X(\m_blake2.m_hash256.m_matrix[10][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(net1177),
    .Q(\m_blake2.m_hash256.m_matrix[10][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1176),
    .A1(\m_blake2.m_hash256.m_matrix[10][23] ),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[10][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][16] ),
    .A1(\m_blake2.m_hash256.m_matrix[10][24] ),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[10][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(net1548),
    .Q(\m_blake2.m_hash256.m_matrix[10][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1547),
    .A1(\m_blake2.m_hash256.m_matrix[10][25] ),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[10][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1711),
    .A1(\m_blake2.m_hash256.m_matrix[10][26] ),
    .S(net607),
    .X(\m_blake2.m_hash256.m_matrix[10][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][19] ),
    .A1(net1266),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[10][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(net1400),
    .Q(\m_blake2.m_hash256.m_matrix[10][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1399),
    .A1(\m_blake2.m_hash256.m_matrix[10][9] ),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[10][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][20] ),
    .A1(net1264),
    .S(net552),
    .X(\m_blake2.m_hash256.m_matrix[10][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1597),
    .A1(\m_blake2.m_hash256.m_matrix[10][29] ),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[10][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(net1380),
    .Q(\m_blake2.m_hash256.m_matrix[10][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1379),
    .A1(\m_blake2.m_hash256.m_matrix[10][30] ),
    .S(net564),
    .X(\m_blake2.m_hash256.m_matrix[10][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1871),
    .A1(\m_blake2.m_hash256.m_matrix[10][31] ),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[10][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][24] ),
    .A1(\m_blake2.m_hash256.m_matrix[11][0] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[10][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(net1257),
    .Q(\m_blake2.m_hash256.m_matrix[10][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][25] ),
    .A1(net1256),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[10][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][26] ),
    .A1(\m_blake2.m_hash256.m_matrix[11][2] ),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[10][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1266),
    .A1(net1216),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[10][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1264),
    .A1(\m_blake2.m_hash256.m_matrix[11][4] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[10][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][29] ),
    .A1(net1675),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[10][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][2] ),
    .A1(net1291),
    .S(net606),
    .X(\m_blake2.m_hash256.m_matrix[10][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(net1057),
    .Q(\m_blake2.m_hash256.m_matrix[10][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][30] ),
    .A1(net1056),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[10][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][31] ),
    .A1(net1698),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[10][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net966),
    .A1(net1265),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[10][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][4] ),
    .A1(net1091),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[10][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][5] ),
    .A1(net1660),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[10][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[10][6] ),
    .A1(net1531),
    .S(net567),
    .X(\m_blake2.m_hash256.m_matrix[10][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1302),
    .A1(net1176),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[10][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1822),
    .A1(\m_blake2.m_hash256.m_matrix[10][16] ),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[10][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[10][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[10][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[10][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[10][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1629),
    .A1(net1547),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[10][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][0] ),
    .A1(\m_blake2.m_hash256.m_matrix[11][8] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[11][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(net1285),
    .Q(\m_blake2.m_hash256.m_matrix[11][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1284),
    .A1(\m_blake2.m_hash256.m_matrix[11][18] ),
    .S(net606),
    .X(\m_blake2.m_hash256.m_matrix[11][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1138),
    .A1(\m_blake2.m_hash256.m_matrix[11][19] ),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[11][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][12] ),
    .A1(net1480),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[11][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][13] ),
    .A1(net1748),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[11][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1248),
    .A1(net1289),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[11][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][15] ),
    .A1(net1858),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[11][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1891),
    .A1(\m_blake2.m_hash256.m_matrix[11][24] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[11][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1368),
    .Q(\m_blake2.m_hash256.m_matrix[11][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1367),
    .A1(\m_blake2.m_hash256.m_matrix[11][25] ),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[11][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(net1158),
    .Q(\m_blake2.m_hash256.m_matrix[11][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][18] ),
    .A1(net1157),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[11][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][19] ),
    .A1(\m_blake2.m_hash256.m_matrix[11][27] ),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[11][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1256),
    .A1(net1341),
    .S(net582),
    .X(\m_blake2.m_hash256.m_matrix[11][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(net1481),
    .Q(\m_blake2.m_hash256.m_matrix[11][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1480),
    .A1(\m_blake2.m_hash256.m_matrix[11][28] ),
    .S(net552),
    .X(\m_blake2.m_hash256.m_matrix[11][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1748),
    .A1(net1624),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[11][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1289),
    .A1(\m_blake2.m_hash256.m_matrix[11][30] ),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[11][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(net1761),
    .Q(\m_blake2.m_hash256.m_matrix[11][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][23] ),
    .A1(net1760),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[11][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][24] ),
    .A1(net1561),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[11][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1806),
    .Q(\m_blake2.m_hash256.m_matrix[11][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][25] ),
    .A1(net1805),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[11][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1157),
    .A1(\m_blake2.m_hash256.m_matrix[12][2] ),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[11][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][27] ),
    .A1(\m_blake2.m_hash256.m_matrix[12][3] ),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[11][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1810),
    .A1(\m_blake2.m_hash256.m_matrix[12][4] ),
    .S(net552),
    .X(\m_blake2.m_hash256.m_matrix[11][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(net1625),
    .Q(\m_blake2.m_hash256.m_matrix[11][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1624),
    .A1(\m_blake2.m_hash256.m_matrix[12][5] ),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[11][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][2] ),
    .A1(net1284),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[11][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][30] ),
    .A1(net1841),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[11][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1760),
    .A1(\m_blake2.m_hash256.m_matrix[12][7] ),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[11][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1216),
    .A1(net1138),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[11][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[11][4] ),
    .A1(\m_blake2.m_hash256.m_matrix[11][12] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[11][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1675),
    .A1(\m_blake2.m_hash256.m_matrix[11][13] ),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[11][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1056),
    .A1(\m_blake2.m_hash256.m_matrix[11][14] ),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[11][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1698),
    .A1(\m_blake2.m_hash256.m_matrix[11][15] ),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[11][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1886),
    .A1(\m_blake2.m_hash256.m_matrix[11][16] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[11][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[11][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[11][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[11][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[11][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1341),
    .A1(net1367),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[11][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1561),
    .A1(net1590),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[12][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net954),
    .A1(net1080),
    .S(net606),
    .X(\m_blake2.m_hash256.m_matrix[12][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1674),
    .A1(\m_blake2.m_hash256.m_matrix[12][19] ),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[12][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][12] ),
    .A1(net1757),
    .S(net552),
    .X(\m_blake2.m_hash256.m_matrix[12][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][13] ),
    .A1(net996),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[12][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][14] ),
    .A1(net1811),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[12][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][15] ),
    .A1(\m_blake2.m_hash256.m_matrix[12][23] ),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[12][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1666),
    .A1(\m_blake2.m_hash256.m_matrix[12][24] ),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1060),
    .Q(\m_blake2.m_hash256.m_matrix[12][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][17] ),
    .A1(net1059),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[12][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1080),
    .A1(net1343),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[12][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][19] ),
    .A1(net1244),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[12][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1739),
    .Q(\m_blake2.m_hash256.m_matrix[12][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][1] ),
    .A1(net1738),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[12][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1757),
    .A1(net1787),
    .S(net552),
    .X(\m_blake2.m_hash256.m_matrix[12][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(net997),
    .Q(\m_blake2.m_hash256.m_matrix[12][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net996),
    .A1(\m_blake2.m_hash256.m_matrix[12][29] ),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[12][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1811),
    .A1(\m_blake2.m_hash256.m_matrix[12][30] ),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[12][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][23] ),
    .A1(net1862),
    .S(net558),
    .X(\m_blake2.m_hash256.m_matrix[12][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][24] ),
    .A1(\m_blake2.m_hash256.m_matrix[13][0] ),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[12][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1059),
    .A1(net1132),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[12][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1343),
    .A1(\m_blake2.m_hash256.m_matrix[13][2] ),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[12][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1244),
    .A1(\m_blake2.m_hash256.m_matrix[13][3] ),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[12][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1787),
    .A1(\m_blake2.m_hash256.m_matrix[13][4] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[12][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(net1129),
    .Q(\m_blake2.m_hash256.m_matrix[12][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1128),
    .A1(\m_blake2.m_hash256.m_matrix[13][5] ),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[12][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][2] ),
    .A1(net954),
    .S(net606),
    .X(\m_blake2.m_hash256.m_matrix[12][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][30] ),
    .A1(net1383),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[12][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1862),
    .A1(net1790),
    .S(net558),
    .X(\m_blake2.m_hash256.m_matrix[12][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1725),
    .A1(net1674),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[12][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1866),
    .A1(\m_blake2.m_hash256.m_matrix[12][12] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[12][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1791),
    .A1(\m_blake2.m_hash256.m_matrix[12][13] ),
    .S(net550),
    .X(\m_blake2.m_hash256.m_matrix[12][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1841),
    .A1(\m_blake2.m_hash256.m_matrix[12][14] ),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[12][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][7] ),
    .A1(\m_blake2.m_hash256.m_matrix[12][15] ),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[12][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[12][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[12][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1590),
    .A1(net1666),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[12][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[12][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1588),
    .Q(\m_blake2.m_hash256.m_matrix[12][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[12][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[12][9] ),
    .A1(net1587),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[12][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][0] ),
    .A1(\m_blake2.m_hash256.m_matrix[13][8] ),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[13][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1832),
    .A1(net1793),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[13][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][11] ),
    .A1(net1664),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[13][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][12] ),
    .A1(\m_blake2.m_hash256.m_matrix[13][20] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[13][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1594),
    .A1(net1506),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[13][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][14] ),
    .A1(net1688),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[13][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][15] ),
    .A1(\m_blake2.m_hash256.m_matrix[13][23] ),
    .S(net558),
    .X(\m_blake2.m_hash256.m_matrix[13][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1511),
    .A1(net1496),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[13][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(net1294),
    .Q(\m_blake2.m_hash256.m_matrix[13][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1293),
    .A1(\m_blake2.m_hash256.m_matrix[13][25] ),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[13][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(net1794),
    .Q(\m_blake2.m_hash256.m_matrix[13][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][18] ),
    .A1(net1734),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[13][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1664),
    .A1(\m_blake2.m_hash256.m_matrix[13][27] ),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[13][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1132),
    .A1(net1421),
    .S(net582),
    .X(\m_blake2.m_hash256.m_matrix[13][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][20] ),
    .A1(net1885),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[13][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1506),
    .A1(net1438),
    .S(net546),
    .X(\m_blake2.m_hash256.m_matrix[13][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1688),
    .A1(\m_blake2.m_hash256.m_matrix[13][30] ),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[13][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][23] ),
    .A1(net1834),
    .S(net558),
    .X(\m_blake2.m_hash256.m_matrix[13][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1496),
    .A1(\m_blake2.m_hash256.m_matrix[14][0] ),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[13][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1752),
    .A1(net1709),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[13][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1734),
    .A1(net1717),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[13][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1671),
    .A1(\m_blake2.m_hash256.m_matrix[14][3] ),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[13][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1885),
    .A1(\m_blake2.m_hash256.m_matrix[14][4] ),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[13][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1438),
    .A1(net1209),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[13][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][2] ),
    .A1(net1832),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[13][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][30] ),
    .A1(net1706),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[13][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1834),
    .A1(\m_blake2.m_hash256.m_matrix[14][7] ),
    .S(net558),
    .X(\m_blake2.m_hash256.m_matrix[13][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][3] ),
    .A1(net1804),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[13][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][4] ),
    .A1(\m_blake2.m_hash256.m_matrix[13][12] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[13][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1646),
    .A1(net1594),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[13][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1383),
    .A1(\m_blake2.m_hash256.m_matrix[13][14] ),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[13][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1790),
    .A1(\m_blake2.m_hash256.m_matrix[13][15] ),
    .S(net550),
    .X(\m_blake2.m_hash256.m_matrix[13][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(net1512),
    .Q(\m_blake2.m_hash256.m_matrix[13][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[13][8] ),
    .A1(net1511),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[13][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[13][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[13][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[13][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1421),
    .A1(net1293),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[13][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][0] ),
    .A1(net1693),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[14][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][10] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][18] ),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[14][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][11] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][19] ),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[14][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][12] ),
    .A1(net1406),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[14][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][13] ),
    .A1(net1700),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[14][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][14] ),
    .A1(net1747),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[14][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][15] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][23] ),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[14][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1765),
    .A1(net1707),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[14][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][17] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][25] ),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[14][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1732),
    .A1(net1165),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[14][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][19] ),
    .A1(net1821),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[14][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1709),
    .A1(\m_blake2.m_hash256.m_matrix[14][9] ),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[14][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1406),
    .A1(net1150),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[14][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1700),
    .A1(\m_blake2.m_hash256.m_matrix[14][29] ),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[14][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1747),
    .A1(\m_blake2.m_hash256.m_matrix[14][30] ),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[14][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][23] ),
    .A1(net1574),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[14][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1707),
    .A1(\m_blake2.m_hash256.m_matrix[15][0] ),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[14][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][25] ),
    .A1(net1799),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[14][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(net1166),
    .Q(\m_blake2.m_hash256.m_matrix[14][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1165),
    .A1(\m_blake2.m_hash256.m_matrix[15][2] ),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1821),
    .A1(\m_blake2.m_hash256.m_matrix[15][3] ),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[14][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1150),
    .A1(\m_blake2.m_hash256.m_matrix[15][4] ),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[14][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][29] ),
    .A1(\m_blake2.m_hash256.m_matrix[15][5] ),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[14][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1717),
    .A1(\m_blake2.m_hash256.m_matrix[14][10] ),
    .S(net604),
    .X(\m_blake2.m_hash256.m_matrix[14][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][30] ),
    .A1(net1502),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[14][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1574),
    .A1(\m_blake2.m_hash256.m_matrix[15][7] ),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[14][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][3] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][11] ),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[14][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][4] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][12] ),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[14][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1209),
    .A1(\m_blake2.m_hash256.m_matrix[14][13] ),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[14][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1706),
    .A1(\m_blake2.m_hash256.m_matrix[14][14] ),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[14][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][7] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][15] ),
    .S(net550),
    .X(\m_blake2.m_hash256.m_matrix[14][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(net1694),
    .Q(\m_blake2.m_hash256.m_matrix[14][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1693),
    .A1(\m_blake2.m_hash256.m_matrix[14][16] ),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[14][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[14][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[14][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[14][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[14][9] ),
    .A1(\m_blake2.m_hash256.m_matrix[14][17] ),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[14][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][0] ),
    .A1(\m_blake2.m_hash256.m_matrix[15][8] ),
    .S(net594),
    .X(\m_blake2.m_hash256.m_matrix[15][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][10] ),
    .A1(\m_blake2.m_hash256.m_matrix[15][18] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][11] ),
    .A1(net1449),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[15][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1355),
    .A1(net1184),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[15][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1475),
    .A1(net1283),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[15][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1836),
    .A1(\m_blake2.m_hash256.m_matrix[15][22] ),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[15][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1641),
    .A1(net1521),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[15][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][16] ),
    .A1(net646),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[15][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1387),
    .A1(net649),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[15][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][18] ),
    .A1(net651),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[15][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(net1450),
    .Q(\m_blake2.m_hash256.m_matrix[15][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1449),
    .A1(\m_blake2.m_hash256.m_matrix[15][27] ),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[15][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1799),
    .A1(\m_blake2.m_hash256.m_matrix[15][9] ),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[15][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1184),
    .A1(\m_blake2.m_hash256.m_matrix[15][28] ),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[15][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1283),
    .A1(\m_blake2.m_hash256.m_matrix[15][29] ),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[15][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][22] ),
    .A1(\m_blake2.m_hash256.m_matrix[15][30] ),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[15][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1521),
    .A1(net935),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[15][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][24] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][25] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][26] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(net643),
    .Q(\m_blake2.m_hash256.m_matrix[15][27] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][28] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][29] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1583),
    .A1(\m_blake2.m_hash256.m_matrix[15][10] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][30] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][31] ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][3] ),
    .A1(\m_blake2.m_hash256.m_matrix[15][11] ),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[15][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][4] ),
    .A1(net1355),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[15][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][5] ),
    .A1(net1475),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[15][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(net1503),
    .Q(\m_blake2.m_hash256.m_matrix[15][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1502),
    .A1(\m_blake2.m_hash256.m_matrix[15][14] ),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[15][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][7] ),
    .A1(net1641),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[15][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][8] ),
    .A1(\m_blake2.m_hash256.m_matrix[15][16] ),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[15][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[15][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[15][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[15][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[15][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[15][9] ),
    .A1(net1387),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[15][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1636),
    .A1(net1500),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(net829),
    .Q(\m_blake2.m_hash256.m_matrix[1][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][10] ),
    .A1(net828),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1407),
    .A1(net1582),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[1][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1070),
    .A1(net1013),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[1][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1520),
    .A1(\m_blake2.m_hash256.m_matrix[1][21] ),
    .S(net546),
    .X(\m_blake2.m_hash256.m_matrix[1][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][14] ),
    .A1(\m_blake2.m_hash256.m_matrix[1][22] ),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[1][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1461),
    .A1(\m_blake2.m_hash256.m_matrix[1][23] ),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[1][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(net1538),
    .Q(\m_blake2.m_hash256.m_matrix[1][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1537),
    .A1(\m_blake2.m_hash256.m_matrix[1][24] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[1][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(net1189),
    .Q(\m_blake2.m_hash256.m_matrix[1][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1188),
    .A1(\m_blake2.m_hash256.m_matrix[1][25] ),
    .S(net556),
    .X(\m_blake2.m_hash256.m_matrix[1][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net828),
    .A1(net1032),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[1][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1582),
    .A1(\m_blake2.m_hash256.m_matrix[1][27] ),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[1][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][1] ),
    .A1(net1328),
    .S(net556),
    .X(\m_blake2.m_hash256.m_matrix[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(net1014),
    .Q(\m_blake2.m_hash256.m_matrix[1][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1013),
    .A1(\m_blake2.m_hash256.m_matrix[1][28] ),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[1][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][21] ),
    .A1(\m_blake2.m_hash256.m_matrix[1][29] ),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[1][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][22] ),
    .A1(\m_blake2.m_hash256.m_matrix[1][30] ),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[1][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][23] ),
    .A1(net1877),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[1][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1723),
    .A1(\m_blake2.m_hash256.m_matrix[2][0] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[1][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1827),
    .A1(net1768),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[1][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1032),
    .A1(net1360),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1392),
    .A1(net1353),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[1][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1603),
    .A1(net1261),
    .S(net560),
    .X(\m_blake2.m_hash256.m_matrix[1][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1837),
    .A1(net1736),
    .S(net546),
    .X(\m_blake2.m_hash256.m_matrix[1][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1612),
    .Q(\m_blake2.m_hash256.m_matrix[1][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1611),
    .A1(\m_blake2.m_hash256.m_matrix[1][10] ),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][30] ),
    .A1(\m_blake2.m_hash256.m_matrix[2][6] ),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[1][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1877),
    .A1(\m_blake2.m_hash256.m_matrix[2][7] ),
    .S(net575),
    .X(\m_blake2.m_hash256.m_matrix[1][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(net1408),
    .Q(\m_blake2.m_hash256.m_matrix[1][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][3] ),
    .A1(net1407),
    .S(net578),
    .X(\m_blake2.m_hash256.m_matrix[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1528),
    .A1(net1070),
    .S(net558),
    .X(\m_blake2.m_hash256.m_matrix[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[1][5] ),
    .A1(net1520),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1676),
    .A1(\m_blake2.m_hash256.m_matrix[1][14] ),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1532),
    .A1(net1461),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(net1501),
    .Q(\m_blake2.m_hash256.m_matrix[1][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1500),
    .A1(\m_blake2.m_hash256.m_matrix[1][16] ),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[1][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[1][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1328),
    .A1(net1188),
    .S(net556),
    .X(\m_blake2.m_hash256.m_matrix[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[2][0] ),
    .A1(net1549),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1340),
    .A1(net1276),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1508),
    .A1(net1446),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[2][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(net1179),
    .Q(\m_blake2.m_hash256.m_matrix[2][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1178),
    .A1(\m_blake2.m_hash256.m_matrix[2][20] ),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[2][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1555),
    .A1(\m_blake2.m_hash256.m_matrix[2][21] ),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[2][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[2][14] ),
    .A1(net1604),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[2][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1552),
    .A1(net1362),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[2][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[2][16] ),
    .A1(net1571),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[2][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(net1485),
    .Q(\m_blake2.m_hash256.m_matrix[2][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1484),
    .A1(\m_blake2.m_hash256.m_matrix[2][25] ),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[2][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1276),
    .A1(net1206),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(net1447),
    .Q(\m_blake2.m_hash256.m_matrix[2][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1446),
    .A1(\m_blake2.m_hash256.m_matrix[2][27] ),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[2][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1768),
    .A1(net1730),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1769),
    .A1(net1905),
    .S(net553),
    .X(\m_blake2.m_hash256.m_matrix[2][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[2][21] ),
    .A1(net1701),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[2][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(net1645),
    .Q(\m_blake2.m_hash256.m_matrix[2][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1604),
    .A1(\m_blake2.m_hash256.m_matrix[2][30] ),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[2][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(net1363),
    .Q(\m_blake2.m_hash256.m_matrix[2][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1362),
    .A1(\m_blake2.m_hash256.m_matrix[2][31] ),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[2][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1571),
    .A1(net1516),
    .S(net598),
    .X(\m_blake2.m_hash256.m_matrix[2][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1731),
    .A1(\m_blake2.m_hash256.m_matrix[3][1] ),
    .S(net556),
    .X(\m_blake2.m_hash256.m_matrix[2][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1206),
    .A1(net1198),
    .S(net589),
    .X(\m_blake2.m_hash256.m_matrix[2][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1605),
    .A1(\m_blake2.m_hash256.m_matrix[3][3] ),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[2][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1864),
    .A1(net1638),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[2][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1701),
    .A1(net1685),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[2][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1360),
    .A1(\m_blake2.m_hash256.m_matrix[2][10] ),
    .S(net605),
    .X(\m_blake2.m_hash256.m_matrix[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(net1840),
    .Q(\m_blake2.m_hash256.m_matrix[2][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1644),
    .A1(\m_blake2.m_hash256.m_matrix[3][6] ),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[2][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1813),
    .A1(net1673),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[2][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(net1354),
    .Q(\m_blake2.m_hash256.m_matrix[2][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1353),
    .A1(\m_blake2.m_hash256.m_matrix[2][11] ),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1261),
    .A1(net1178),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1736),
    .A1(net1555),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1894),
    .A1(\m_blake2.m_hash256.m_matrix[2][14] ),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1887),
    .A1(net1552),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1549),
    .A1(\m_blake2.m_hash256.m_matrix[2][16] ),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[2][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[2][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1730),
    .A1(net1484),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(net1517),
    .Q(\m_blake2.m_hash256.m_matrix[3][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1516),
    .A1(\m_blake2.m_hash256.m_matrix[3][8] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[3][10] ),
    .A1(net1401),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[3][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1640),
    .A1(net1589),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[3][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1572),
    .A1(\m_blake2.m_hash256.m_matrix[3][20] ),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[3][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1661),
    .A1(net1610),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[3][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[3][14] ),
    .A1(net1635),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[3][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1650),
    .A1(net1126),
    .S(net567),
    .X(\m_blake2.m_hash256.m_matrix[3][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1667),
    .A1(net1559),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1692),
    .A1(\m_blake2.m_hash256.m_matrix[3][25] ),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[3][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1401),
    .A1(net1333),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[3][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1589),
    .A1(net1364),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[3][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1789),
    .Q(\m_blake2.m_hash256.m_matrix[3][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1788),
    .A1(\m_blake2.m_hash256.m_matrix[3][9] ),
    .S(net582),
    .X(\m_blake2.m_hash256.m_matrix[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[3][20] ),
    .A1(net1397),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[3][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1610),
    .A1(net1592),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[3][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1635),
    .A1(net1637),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[3][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1126),
    .A1(net1035),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[3][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(net1560),
    .Q(\m_blake2.m_hash256.m_matrix[3][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1559),
    .A1(\m_blake2.m_hash256.m_matrix[4][0] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[3][25] ),
    .A1(net1786),
    .S(net581),
    .X(\m_blake2.m_hash256.m_matrix[3][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1334),
    .Q(\m_blake2.m_hash256.m_matrix[3][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1333),
    .A1(\m_blake2.m_hash256.m_matrix[4][2] ),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[3][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1364),
    .A1(\m_blake2.m_hash256.m_matrix[4][3] ),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[3][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1397),
    .A1(\m_blake2.m_hash256.m_matrix[4][4] ),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[3][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1592),
    .A1(net1518),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[3][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1198),
    .A1(\m_blake2.m_hash256.m_matrix[3][10] ),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1637),
    .A1(net1619),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[3][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1035),
    .A1(\m_blake2.m_hash256.m_matrix[4][7] ),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[3][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1695),
    .A1(net1640),
    .S(net602),
    .X(\m_blake2.m_hash256.m_matrix[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1638),
    .A1(net1572),
    .S(net557),
    .X(\m_blake2.m_hash256.m_matrix[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1685),
    .A1(\m_blake2.m_hash256.m_matrix[3][13] ),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1839),
    .A1(\m_blake2.m_hash256.m_matrix[3][14] ),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1673),
    .A1(net1650),
    .S(net579),
    .X(\m_blake2.m_hash256.m_matrix[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1784),
    .A1(\m_blake2.m_hash256.m_matrix[3][16] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[3][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[3][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1833),
    .A1(net1692),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1828),
    .A1(net1623),
    .S(net590),
    .X(\m_blake2.m_hash256.m_matrix[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1474),
    .A1(net1259),
    .S(net602),
    .X(\m_blake2.m_hash256.m_matrix[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[4][11] ),
    .A1(\m_blake2.m_hash256.m_matrix[4][19] ),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[4][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1743),
    .A1(net1714),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[4][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1713),
    .A1(net1581),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[4][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1716),
    .A1(net1651),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[4][15] ),
    .A1(net1255),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[4][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1602),
    .A1(net1593),
    .S(net584),
    .X(\m_blake2.m_hash256.m_matrix[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1729),
    .A1(\m_blake2.m_hash256.m_matrix[4][25] ),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[4][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1260),
    .Q(\m_blake2.m_hash256.m_matrix[4][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1259),
    .A1(\m_blake2.m_hash256.m_matrix[4][26] ),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[4][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[4][19] ),
    .A1(net1171),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[4][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1786),
    .A1(\m_blake2.m_hash256.m_matrix[4][9] ),
    .S(net581),
    .X(\m_blake2.m_hash256.m_matrix[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1714),
    .A1(net1535),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[4][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1581),
    .A1(net1568),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[4][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1651),
    .A1(net1578),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[4][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1255),
    .A1(\m_blake2.m_hash256.m_matrix[4][31] ),
    .S(net575),
    .X(\m_blake2.m_hash256.m_matrix[4][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1593),
    .A1(net1433),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[4][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(net1751),
    .Q(\m_blake2.m_hash256.m_matrix[4][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1750),
    .A1(\m_blake2.m_hash256.m_matrix[5][1] ),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[4][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1304),
    .Q(\m_blake2.m_hash256.m_matrix[4][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1303),
    .A1(\m_blake2.m_hash256.m_matrix[5][2] ),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[4][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1172),
    .Q(\m_blake2.m_hash256.m_matrix[4][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1171),
    .A1(\m_blake2.m_hash256.m_matrix[5][3] ),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[4][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1535),
    .A1(net1525),
    .S(net553),
    .X(\m_blake2.m_hash256.m_matrix[4][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1568),
    .A1(net1050),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[4][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1498),
    .A1(net1474),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1578),
    .A1(net1488),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[4][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[4][31] ),
    .A1(net1715),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[4][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1888),
    .A1(\m_blake2.m_hash256.m_matrix[4][11] ),
    .S(net602),
    .X(\m_blake2.m_hash256.m_matrix[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[4][4] ),
    .A1(net1743),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(net1519),
    .Q(\m_blake2.m_hash256.m_matrix[4][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1518),
    .A1(\m_blake2.m_hash256.m_matrix[4][13] ),
    .S(net547),
    .X(\m_blake2.m_hash256.m_matrix[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(net1620),
    .Q(\m_blake2.m_hash256.m_matrix[4][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1619),
    .A1(\m_blake2.m_hash256.m_matrix[4][14] ),
    .S(net569),
    .X(\m_blake2.m_hash256.m_matrix[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[4][7] ),
    .A1(\m_blake2.m_hash256.m_matrix[4][15] ),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1623),
    .A1(net1602),
    .S(net584),
    .X(\m_blake2.m_hash256.m_matrix[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[4][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[4][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[4][9] ),
    .A1(net1729),
    .S(net554),
    .X(\m_blake2.m_hash256.m_matrix[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1433),
    .A1(net1217),
    .S(net584),
    .X(\m_blake2.m_hash256.m_matrix[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1566),
    .A1(net1384),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[5][11] ),
    .A1(net1533),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[5][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1403),
    .A1(net1335),
    .S(net553),
    .X(\m_blake2.m_hash256.m_matrix[5][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net963),
    .A1(\m_blake2.m_hash256.m_matrix[5][21] ),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[5][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1705),
    .A1(net1655),
    .S(net570),
    .X(\m_blake2.m_hash256.m_matrix[5][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[5][15] ),
    .A1(net1371),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[5][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1429),
    .A1(net1325),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(net1819),
    .Q(\m_blake2.m_hash256.m_matrix[5][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1818),
    .A1(\m_blake2.m_hash256.m_matrix[5][25] ),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[5][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1384),
    .A1(net1273),
    .S(net589),
    .X(\m_blake2.m_hash256.m_matrix[5][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(net1534),
    .Q(\m_blake2.m_hash256.m_matrix[5][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1533),
    .A1(\m_blake2.m_hash256.m_matrix[5][27] ),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[5][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1857),
    .A1(net1846),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(net1336),
    .Q(\m_blake2.m_hash256.m_matrix[5][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1335),
    .A1(\m_blake2.m_hash256.m_matrix[5][28] ),
    .S(net553),
    .X(\m_blake2.m_hash256.m_matrix[5][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[5][21] ),
    .A1(net1553),
    .S(net548),
    .X(\m_blake2.m_hash256.m_matrix[5][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1655),
    .A1(\m_blake2.m_hash256.m_matrix[5][30] ),
    .S(net570),
    .X(\m_blake2.m_hash256.m_matrix[5][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1371),
    .A1(net1049),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[5][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1326),
    .Q(\m_blake2.m_hash256.m_matrix[5][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1325),
    .A1(\m_blake2.m_hash256.m_matrix[6][0] ),
    .S(net585),
    .X(\m_blake2.m_hash256.m_matrix[5][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(net1884),
    .Q(\m_blake2.m_hash256.m_matrix[5][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1883),
    .A1(\m_blake2.m_hash256.m_matrix[6][1] ),
    .S(net581),
    .X(\m_blake2.m_hash256.m_matrix[5][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1274),
    .Q(\m_blake2.m_hash256.m_matrix[5][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1273),
    .A1(\m_blake2.m_hash256.m_matrix[6][2] ),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[5][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1830),
    .A1(net1746),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[5][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1413),
    .A1(\m_blake2.m_hash256.m_matrix[6][4] ),
    .S(net553),
    .X(\m_blake2.m_hash256.m_matrix[5][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(net1554),
    .Q(\m_blake2.m_hash256.m_matrix[5][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1553),
    .A1(\m_blake2.m_hash256.m_matrix[6][5] ),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[5][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1609),
    .A1(net1566),
    .S(net601),
    .X(\m_blake2.m_hash256.m_matrix[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1720),
    .A1(\m_blake2.m_hash256.m_matrix[6][6] ),
    .S(net564),
    .X(\m_blake2.m_hash256.m_matrix[5][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1049),
    .A1(\m_blake2.m_hash256.m_matrix[6][7] ),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[5][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1812),
    .A1(\m_blake2.m_hash256.m_matrix[5][11] ),
    .S(net559),
    .X(\m_blake2.m_hash256.m_matrix[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_4_clk),
    .D(net1526),
    .Q(\m_blake2.m_hash256.m_matrix[5][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1525),
    .A1(\m_blake2.m_hash256.m_matrix[5][12] ),
    .S(net553),
    .X(\m_blake2.m_hash256.m_matrix[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1050),
    .A1(net963),
    .S(net542),
    .X(\m_blake2.m_hash256.m_matrix[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(net1489),
    .Q(\m_blake2.m_hash256.m_matrix[5][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1488),
    .A1(\m_blake2.m_hash256.m_matrix[5][14] ),
    .S(net568),
    .X(\m_blake2.m_hash256.m_matrix[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1715),
    .A1(\m_blake2.m_hash256.m_matrix[5][15] ),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1217),
    .A1(net1904),
    .S(net584),
    .X(\m_blake2.m_hash256.m_matrix[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[5][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[5][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1846),
    .A1(net1818),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1417),
    .Q(\m_blake2.m_hash256.m_matrix[6][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1416),
    .A1(\m_blake2.m_hash256.m_matrix[6][8] ),
    .S(net590),
    .X(\m_blake2.m_hash256.m_matrix[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][10] ),
    .A1(net1564),
    .S(net589),
    .X(\m_blake2.m_hash256.m_matrix[6][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1728),
    .A1(net1357),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[6][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1418),
    .A1(\m_blake2.m_hash256.m_matrix[6][20] ),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[6][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1186),
    .A1(net1148),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[6][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1719),
    .A1(\m_blake2.m_hash256.m_matrix[6][22] ),
    .S(net564),
    .X(\m_blake2.m_hash256.m_matrix[6][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][15] ),
    .A1(\m_blake2.m_hash256.m_matrix[6][23] ),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[6][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1844),
    .A1(\m_blake2.m_hash256.m_matrix[6][24] ),
    .S(net595),
    .X(\m_blake2.m_hash256.m_matrix[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][17] ),
    .A1(net1668),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[6][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1564),
    .A1(net1546),
    .S(net597),
    .X(\m_blake2.m_hash256.m_matrix[6][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(net1358),
    .Q(\m_blake2.m_hash256.m_matrix[6][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1357),
    .A1(\m_blake2.m_hash256.m_matrix[6][27] ),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[6][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(net1756),
    .Q(\m_blake2.m_hash256.m_matrix[6][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][1] ),
    .A1(net1755),
    .S(net581),
    .X(\m_blake2.m_hash256.m_matrix[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][20] ),
    .A1(net1686),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[6][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1148),
    .A1(\m_blake2.m_hash256.m_matrix[6][29] ),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[6][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][22] ),
    .A1(net981),
    .S(net570),
    .X(\m_blake2.m_hash256.m_matrix[6][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1878),
    .A1(\m_blake2.m_hash256.m_matrix[6][31] ),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[6][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][24] ),
    .A1(net1236),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[6][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_5_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1668),
    .A1(\m_blake2.m_hash256.m_matrix[7][1] ),
    .S(net555),
    .X(\m_blake2.m_hash256.m_matrix[6][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1546),
    .A1(net1455),
    .S(net597),
    .X(\m_blake2.m_hash256.m_matrix[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1628),
    .Q(\m_blake2.m_hash256.m_matrix[6][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1627),
    .A1(\m_blake2.m_hash256.m_matrix[7][3] ),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[6][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1686),
    .A1(net1569),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[6][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][29] ),
    .A1(net1781),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[6][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1565),
    .A1(\m_blake2.m_hash256.m_matrix[6][10] ),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net981),
    .A1(\m_blake2.m_hash256.m_matrix[7][6] ),
    .S(net570),
    .X(\m_blake2.m_hash256.m_matrix[6][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][31] ),
    .A1(\m_blake2.m_hash256.m_matrix[7][7] ),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[6][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1746),
    .A1(net1728),
    .S(net573),
    .X(\m_blake2.m_hash256.m_matrix[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][4] ),
    .A1(net1418),
    .S(net549),
    .X(\m_blake2.m_hash256.m_matrix[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(net1187),
    .Q(\m_blake2.m_hash256.m_matrix[6][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][5] ),
    .A1(net1186),
    .S(net546),
    .X(\m_blake2.m_hash256.m_matrix[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][6] ),
    .A1(net1719),
    .S(net570),
    .X(\m_blake2.m_hash256.m_matrix[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[6][7] ),
    .A1(\m_blake2.m_hash256.m_matrix[6][15] ),
    .S(net577),
    .X(\m_blake2.m_hash256.m_matrix[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1873),
    .A1(net1844),
    .S(net584),
    .X(\m_blake2.m_hash256.m_matrix[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[6][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[6][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1755),
    .A1(\m_blake2.m_hash256.m_matrix[6][17] ),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(net1237),
    .Q(\m_blake2.m_hash256.m_matrix[7][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1236),
    .A1(\m_blake2.m_hash256.m_matrix[7][8] ),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][10] ),
    .A1(\m_blake2.m_hash256.m_matrix[7][18] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1393),
    .A1(net1155),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[7][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(net1616),
    .Q(\m_blake2.m_hash256.m_matrix[7][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1615),
    .A1(\m_blake2.m_hash256.m_matrix[7][20] ),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[7][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][13] ),
    .A1(net1680),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[7][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1415),
    .A1(\m_blake2.m_hash256.m_matrix[7][22] ),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[7][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1201),
    .A1(\m_blake2.m_hash256.m_matrix[7][23] ),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[7][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1691),
    .A1(\m_blake2.m_hash256.m_matrix[7][24] ),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1633),
    .A1(\m_blake2.m_hash256.m_matrix[7][25] ),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[7][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][18] ),
    .A1(net1241),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[7][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(net1156),
    .Q(\m_blake2.m_hash256.m_matrix[7][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1155),
    .A1(\m_blake2.m_hash256.m_matrix[7][27] ),
    .S(net602),
    .X(\m_blake2.m_hash256.m_matrix[7][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1835),
    .A1(\m_blake2.m_hash256.m_matrix[7][9] ),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(net1663),
    .Q(\m_blake2.m_hash256.m_matrix[7][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1662),
    .A1(\m_blake2.m_hash256.m_matrix[7][28] ),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[7][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1680),
    .A1(\m_blake2.m_hash256.m_matrix[7][29] ),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[7][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1708),
    .A1(net1558),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[7][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][23] ),
    .A1(net1297),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[7][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][24] ),
    .A1(net1766),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[7][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][25] ),
    .A1(\m_blake2.m_hash256.m_matrix[8][1] ),
    .S(net587),
    .X(\m_blake2.m_hash256.m_matrix[7][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(net1242),
    .Q(\m_blake2.m_hash256.m_matrix[7][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1241),
    .A1(\m_blake2.m_hash256.m_matrix[8][2] ),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[7][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1456),
    .A1(net1174),
    .S(net602),
    .X(\m_blake2.m_hash256.m_matrix[7][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1843),
    .A1(\m_blake2.m_hash256.m_matrix[8][4] ),
    .S(net544),
    .X(\m_blake2.m_hash256.m_matrix[7][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][29] ),
    .A1(\m_blake2.m_hash256.m_matrix[8][5] ),
    .S(net541),
    .X(\m_blake2.m_hash256.m_matrix[7][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1455),
    .A1(\m_blake2.m_hash256.m_matrix[7][10] ),
    .S(net597),
    .X(\m_blake2.m_hash256.m_matrix[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1558),
    .A1(net1524),
    .S(net567),
    .X(\m_blake2.m_hash256.m_matrix[7][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1297),
    .A1(net1269),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[7][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1642),
    .A1(net1393),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(net1570),
    .Q(\m_blake2.m_hash256.m_matrix[7][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1569),
    .A1(\m_blake2.m_hash256.m_matrix[7][12] ),
    .S(net545),
    .X(\m_blake2.m_hash256.m_matrix[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1781),
    .A1(\m_blake2.m_hash256.m_matrix[7][13] ),
    .S(net541),
    .X(\m_blake2.m_hash256.m_matrix[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][6] ),
    .A1(net1415),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][7] ),
    .A1(net1201),
    .S(net571),
    .X(\m_blake2.m_hash256.m_matrix[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(net1580),
    .Q(\m_blake2.m_hash256.m_matrix[7][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1579),
    .A1(\m_blake2.m_hash256.m_matrix[7][16] ),
    .S(net592),
    .X(\m_blake2.m_hash256.m_matrix[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[7][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(\m_blake2.m_hash256.m_matrix[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[7][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[7][9] ),
    .A1(net1633),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(net1767),
    .Q(\m_blake2.m_hash256.m_matrix[8][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1766),
    .A1(\m_blake2.m_hash256.m_matrix[8][8] ),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][10] ),
    .A1(\m_blake2.m_hash256.m_matrix[8][18] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_6_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1630),
    .A1(net1618),
    .S(net574),
    .X(\m_blake2.m_hash256.m_matrix[8][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][12] ),
    .A1(net1771),
    .S(net544),
    .X(\m_blake2.m_hash256.m_matrix[8][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(net1043),
    .Q(\m_blake2.m_hash256.m_matrix[8][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][13] ),
    .A1(net1042),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[8][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(net1200),
    .Q(\m_blake2.m_hash256.m_matrix[8][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][14] ),
    .A1(net1199),
    .S(net563),
    .X(\m_blake2.m_hash256.m_matrix[8][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1585),
    .A1(\m_blake2.m_hash256.m_matrix[8][23] ),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[8][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(net1483),
    .Q(\m_blake2.m_hash256.m_matrix[8][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][16] ),
    .A1(net1482),
    .S(net594),
    .X(\m_blake2.m_hash256.m_matrix[8][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(net1282),
    .Q(\m_blake2.m_hash256.m_matrix[8][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1281),
    .A1(\m_blake2.m_hash256.m_matrix[8][25] ),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[8][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][18] ),
    .A1(net1212),
    .S(net597),
    .X(\m_blake2.m_hash256.m_matrix[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1618),
    .A1(net1425),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[8][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][1] ),
    .A1(\m_blake2.m_hash256.m_matrix[8][9] ),
    .S(net586),
    .X(\m_blake2.m_hash256.m_matrix[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1771),
    .A1(net1758),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[8][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1042),
    .A1(\m_blake2.m_hash256.m_matrix[8][29] ),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[8][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_73_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1199),
    .A1(\m_blake2.m_hash256.m_matrix[8][30] ),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[8][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][23] ),
    .A1(net1193),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[8][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1482),
    .A1(\m_blake2.m_hash256.m_matrix[9][0] ),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[8][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(net1332),
    .Q(\m_blake2.m_hash256.m_matrix[8][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][25] ),
    .A1(net1331),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[8][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_17_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1212),
    .A1(\m_blake2.m_hash256.m_matrix[9][2] ),
    .S(net597),
    .X(\m_blake2.m_hash256.m_matrix[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][27] ),
    .A1(net1224),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[8][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(net1759),
    .Q(\m_blake2.m_hash256.m_matrix[8][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1758),
    .A1(\m_blake2.m_hash256.m_matrix[9][4] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[8][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_74_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][29] ),
    .A1(\m_blake2.m_hash256.m_matrix[9][5] ),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[8][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1814),
    .A1(\m_blake2.m_hash256.m_matrix[8][10] ),
    .S(net596),
    .X(\m_blake2.m_hash256.m_matrix[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1337),
    .A1(net1684),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[8][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(net1194),
    .Q(\m_blake2.m_hash256.m_matrix[8][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1193),
    .A1(\m_blake2.m_hash256.m_matrix[9][7] ),
    .S(net572),
    .X(\m_blake2.m_hash256.m_matrix[8][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_13_clk),
    .D(net1175),
    .Q(\m_blake2.m_hash256.m_matrix[8][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1174),
    .A1(\m_blake2.m_hash256.m_matrix[8][11] ),
    .S(net600),
    .X(\m_blake2.m_hash256.m_matrix[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1901),
    .A1(\m_blake2.m_hash256.m_matrix[8][12] ),
    .S(net544),
    .X(\m_blake2.m_hash256.m_matrix[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(net1492),
    .Q(\m_blake2.m_hash256.m_matrix[8][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][5] ),
    .A1(net1491),
    .S(net541),
    .X(\m_blake2.m_hash256.m_matrix[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1524),
    .A1(\m_blake2.m_hash256.m_matrix[8][14] ),
    .S(net565),
    .X(\m_blake2.m_hash256.m_matrix[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_71_clk),
    .D(net1270),
    .Q(\m_blake2.m_hash256.m_matrix[8][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1269),
    .A1(\m_blake2.m_hash256.m_matrix[8][15] ),
    .S(net566),
    .X(\m_blake2.m_hash256.m_matrix[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_18_clk),
    .D(net1703),
    .Q(\m_blake2.m_hash256.m_matrix[8][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[8][8] ),
    .A1(net1702),
    .S(net593),
    .X(\m_blake2.m_hash256.m_matrix[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[8][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_16_clk),
    .D(\m_blake2.m_hash256.m_matrix[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[8][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1374),
    .A1(net1281),
    .S(net588),
    .X(\m_blake2.m_hash256.m_matrix[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][0] ),
    .A1(net1775),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1850),
    .A1(net1848),
    .S(net606),
    .X(\m_blake2.m_hash256.m_matrix[9][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(net1477),
    .Q(\m_blake2.m_hash256.m_matrix[9][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1476),
    .A1(\m_blake2.m_hash256.m_matrix[9][19] ),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[9][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1515),
    .A1(net1452),
    .S(net544),
    .X(\m_blake2.m_hash256.m_matrix[9][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(net1808),
    .Q(\m_blake2.m_hash256.m_matrix[9][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1807),
    .A1(\m_blake2.m_hash256.m_matrix[9][21] ),
    .S(net541),
    .X(\m_blake2.m_hash256.m_matrix[9][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][14] ),
    .A1(net1419),
    .S(net564),
    .X(\m_blake2.m_hash256.m_matrix[9][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1315),
    .A1(net1220),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[9][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1782),
    .A1(\m_blake2.m_hash256.m_matrix[9][24] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[9][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net988),
    .A1(net1004),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[9][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1848),
    .A1(\m_blake2.m_hash256.m_matrix[9][26] ),
    .S(net607),
    .X(\m_blake2.m_hash256.m_matrix[9][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1573),
    .A1(\m_blake2.m_hash256.m_matrix[9][27] ),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[9][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1331),
    .A1(\m_blake2.m_hash256.m_matrix[9][9] ),
    .S(net581),
    .X(\m_blake2.m_hash256.m_matrix[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_1_clk),
    .D(net1453),
    .Q(\m_blake2.m_hash256.m_matrix[9][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1452),
    .A1(\m_blake2.m_hash256.m_matrix[9][28] ),
    .S(net543),
    .X(\m_blake2.m_hash256.m_matrix[9][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1823),
    .A1(\m_blake2.m_hash256.m_matrix[9][29] ),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[9][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(net1420),
    .Q(\m_blake2.m_hash256.m_matrix[9][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1419),
    .A1(\m_blake2.m_hash256.m_matrix[9][30] ),
    .S(net564),
    .X(\m_blake2.m_hash256.m_matrix[9][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(net1221),
    .Q(\m_blake2.m_hash256.m_matrix[9][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1220),
    .A1(\m_blake2.m_hash256.m_matrix[9][31] ),
    .S(net575),
    .X(\m_blake2.m_hash256.m_matrix[9][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][24] ),
    .A1(net1802),
    .S(net594),
    .X(\m_blake2.m_hash256.m_matrix[9][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_15_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1004),
    .A1(net1399),
    .S(net583),
    .X(\m_blake2.m_hash256.m_matrix[9][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][26] ),
    .A1(\m_blake2.m_hash256.m_matrix[10][2] ),
    .S(net607),
    .X(\m_blake2.m_hash256.m_matrix[9][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_12_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][27] ),
    .A1(net966),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[9][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1831),
    .A1(\m_blake2.m_hash256.m_matrix[10][4] ),
    .S(net544),
    .X(\m_blake2.m_hash256.m_matrix[9][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][29] ),
    .A1(\m_blake2.m_hash256.m_matrix[10][5] ),
    .S(net541),
    .X(\m_blake2.m_hash256.m_matrix[9][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][2] ),
    .A1(\m_blake2.m_hash256.m_matrix[9][10] ),
    .S(net606),
    .X(\m_blake2.m_hash256.m_matrix[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1754),
    .A1(\m_blake2.m_hash256.m_matrix[10][6] ),
    .S(net564),
    .X(\m_blake2.m_hash256.m_matrix[9][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_2_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1385),
    .A1(net1302),
    .S(net575),
    .X(\m_blake2.m_hash256.m_matrix[9][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(net1225),
    .Q(\m_blake2.m_hash256.m_matrix[9][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1224),
    .A1(\m_blake2.m_hash256.m_matrix[9][11] ),
    .S(net603),
    .X(\m_blake2.m_hash256.m_matrix[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_3_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1800),
    .A1(\m_blake2.m_hash256.m_matrix[9][12] ),
    .S(net551),
    .X(\m_blake2.m_hash256.m_matrix[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_0_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][5] ),
    .A1(net1807),
    .S(net540),
    .X(\m_blake2.m_hash256.m_matrix[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_72_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1684),
    .A1(\m_blake2.m_hash256.m_matrix[9][14] ),
    .S(net562),
    .X(\m_blake2.m_hash256.m_matrix[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_7_clk),
    .D(\m_blake2.m_hash256.m_matrix[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.m_matrix[9][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1382),
    .A1(net1315),
    .S(net576),
    .X(\m_blake2.m_hash256.m_matrix[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(net1776),
    .Q(\m_blake2.m_hash256.m_matrix[9][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1775),
    .A1(\m_blake2.m_hash256.m_matrix[9][16] ),
    .S(net591),
    .X(\m_blake2.m_hash256.m_matrix[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.m_matrix[9][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_14_clk),
    .D(net989),
    .Q(\m_blake2.m_hash256.m_matrix[9][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.m_matrix[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_matrix[9][9] ),
    .A1(net988),
    .S(net580),
    .X(\m_blake2.m_hash256.m_matrix[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.res_cnt_q[0] ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X  (.A(net478),
    .B(\m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__xor2_2_B  (.A(net446),
    .B(\m_blake2.m_hash256.res_cnt_q[0] ),
    .X(\m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__a21oi_2_B1  (.A1(net446),
    .A2(\m_blake2.m_hash256.res_cnt_q[0] ),
    .B1(\m_blake2.m_hash256.res_cnt_q[1] ),
    .Y(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__and3_2_C_X ),
    .B(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__and3_2_C  (.A(net446),
    .B(\m_blake2.m_hash256.res_cnt_q[0] ),
    .C(\m_blake2.m_hash256.res_cnt_q[1] ),
    .X(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.res_cnt_q[1] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__inv_2_Y  (.A(net478),
    .Y(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A  (.A(\m_blake2.m_hash256.res_cnt_q[2] ),
    .B(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__and3_2_C_X ),
    .X(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.res_cnt_q[2] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.res_cnt_q[2] ),
    .B(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__and3_2_C_X ),
    .Y(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .B(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.res_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.res_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.res_cnt_q[3] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.res_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_blake2.m_hash256.res_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.res_cnt_q[3] ),
    .A2(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .B1(\m_blake2.m_hash256.res_cnt_q[4] ),
    .Y(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__and3_2_B_X ),
    .B(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .X(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_io.m_config.nn_q[4] ),
    .B(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A_C ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_io.m_config.nn_q[4] ),
    .B(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__and3_2_B  (.A(\m_blake2.m_hash256.res_cnt_q[3] ),
    .B(\m_blake2.m_hash256.res_cnt_q[4] ),
    .C(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.res_cnt_q[4] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.res_cnt_q[5] ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__xnor2_2_A  (.A(net1689),
    .B(\m_blake2.m_hash256.res_cnt_q[4]_sky130_fd_sc_hd__and3_2_B_X ),
    .Y(\m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__and2b_2_B  (.A_N(net466),
    .B(net462),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[0] ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a21bo_2_X  (.A1(net1815),
    .A2(net152),
    .B1_N(net482),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2b_4 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B  (.A_N(net466),
    .B(net462),
    .Y(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1  (.A1(net462),
    .A2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X ),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_1  (.A1(net462),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .C(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .D(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1_X ),
    .A2(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X ),
    .B1(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_B1_sky130_fd_sc_hd__or3_2_X  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .C(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or4_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_B1 ));
 sky130_fd_sc_hd__o21ai_2 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2  (.A1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1_X ),
    .A2(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X ),
    .B1(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_B1 ),
    .Y(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1  (.A1(net462),
    .A2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1  (.A1(\m_blake2.m_hash256.round_q[0] ),
    .A2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_B  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1_X ),
    .C(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .D(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_B_X ));
 sky130_fd_sc_hd__nor4_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B  (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_A ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X ),
    .C(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_1_X ),
    .D(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_D ),
    .Y(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_A_sky130_fd_sc_hd__o21a_2_X  (.A1(net455),
    .A2(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_A ));
 sky130_fd_sc_hd__o311a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_D_sky130_fd_sc_hd__o311a_2_X  (.A1(net459),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .A3(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(net401),
    .C1(net468),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B  (.A(net456),
    .B(\m_blake2.m_hash256.round_q[0] ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C  (.A(net458),
    .B(net459),
    .C(net462),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X ),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3  (.A1(net451),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .A3(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X ),
    .B1(net444),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B  (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_A ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .C(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_C ),
    .Y(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_A_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .A2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_A ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_C_sky130_fd_sc_hd__o31a_2_X  (.A1(net407),
    .A2(net460),
    .A3(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[1] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net462),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net482),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(net461),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__o311a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1  (.A1(net461),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ),
    .A3(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(net401),
    .C1(net468),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B  (.A(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X ),
    .C(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D_sky130_fd_sc_hd__o31a_2_X  (.A1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1  (.A1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X ),
    .B2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1  (.A1(net461),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .A3(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X ));
 sky130_fd_sc_hd__nor3b_4 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__nor3b_2_Y  (.A(net466),
    .B(net474),
    .C_N(net470),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ));
 sky130_fd_sc_hd__or2_4 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_B2_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2  (.A1(net458),
    .A2(net461),
    .A3(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_X ));
 sky130_fd_sc_hd__nand2_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1 ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net468),
    .B(net474),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1 ));
 sky130_fd_sc_hd__o41a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__o41a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A2(net451),
    .A3(net456),
    .A4(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_D ));
 sky130_fd_sc_hd__o41a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3  (.A1(net453),
    .A2(net457),
    .A3(net461),
    .A4(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1 ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X ));
 sky130_fd_sc_hd__o41a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_1  (.A1(net453),
    .A2(net457),
    .A3(net461),
    .A4(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_1_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_B  (.A(net445),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1 ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net471),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__or2_2_X  (.A(net467),
    .B(net475),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B  (.A(net444),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1 ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C  (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X ),
    .C(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_2  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_2_X ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_3  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_3_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C  (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X ),
    .C(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ));
 sky130_fd_sc_hd__and4_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.round_q[1] ),
    .B(net462),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B  (.A(net460),
    .B(net461),
    .C(\m_blake2.m_hash256.round_q[0] ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o211a_2_A2  (.A1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(net468),
    .C1(net401),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o211a_2_A2_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(net452),
    .A2(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C  (.A(net455),
    .B(net459),
    .C(net461),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .C(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1  (.A1(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_Y ),
    .A2(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_Y ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__a21oi_2 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_Y ),
    .A2(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_Y ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .Y(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[2] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.round_q[1] ),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net482),
    .X(\m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(net459),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[3] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net459),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net482),
    .X(\m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(net457),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[4] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net458),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net482),
    .X(\m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(net456),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[5] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net456),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net482),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.round_q[5] ),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1  (.A1(net454),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__a311o_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1  (.A1(net468),
    .A2(net401),
    .A3(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X ),
    .B1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .C1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_X ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1  (.A1(net454),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_1  (.A1(net454),
    .A2(net456),
    .A3(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C  (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o21a_2_A1_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X ),
    .D(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_D ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X ));
 sky130_fd_sc_hd__o311a_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_D_sky130_fd_sc_hd__o311a_2_X  (.A1(net455),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(net401),
    .C1(net468),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X ),
    .Y(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__nand4_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nand4_2_C  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nand4_2_C_Y ));
 sky130_fd_sc_hd__o41a_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2  (.A1(net451),
    .A2(net454),
    .A3(net460),
    .A4(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_X ));
 sky130_fd_sc_hd__and3b_2 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1_sky130_fd_sc_hd__and3b_2_X  (.A_N(net470),
    .B(net474),
    .C(net466),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B  (.A(net452),
    .B(net454),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A  (.A(net454),
    .B(net456),
    .C(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net444),
    .A2(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .B2(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__o31a_2_A3  (.A1(net452),
    .A2(net458),
    .A3(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or4_2_A  (.A(net454),
    .B(net457),
    .C(net459),
    .D(net461),
    .X(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(net1045),
    .Q(\m_blake2.m_hash256.round_q[6] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1044),
    .A2(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B1(\m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(\m_blake2.m_hash256.fsm_q[2] ),
    .X(\m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(net451),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[7] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net452),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net482),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(net450),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1  (.A1(\m_blake2.m_hash256.round_q[7] ),
    .A2(net451),
    .A3(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(net444),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D  (.A(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .B(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_B ),
    .C(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .D(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .A2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_B ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D  (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_A ),
    .B(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_B ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C ),
    .D(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_A_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ),
    .A2(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_A ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_B_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_B ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X  (.A1(net468),
    .A2(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A ),
    .A3(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_B1 ),
    .B2(net401),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__or2_2_X  (.A(net451),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__or3b_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_B1_sky130_fd_sc_hd__or3b_2_X  (.A(net458),
    .B(net460),
    .C_N(net468),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_B1 ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1  (.A1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A  (.A(net450),
    .B(\m_blake2.m_hash256.round_q[1] ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A  (.A(net450),
    .B(net457),
    .C(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__or3_2 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1  (.A(net450),
    .B(net456),
    .C(net462),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a221o_2_B1  (.A1(net444),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X ),
    .B1(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X ),
    .B2(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .C1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_1_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a221o_2_B1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A  (.A(net450),
    .B(net453),
    .C(net455),
    .D(net457),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1  (.A(net450),
    .B(net456),
    .C(net457),
    .D(net460),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C  (.A(net407),
    .B(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__nor3_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C  (.A(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .Y(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2_X ));
 sky130_fd_sc_hd__and4_2 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__a21o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o21ai_2_A2_Y ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C  (.A(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or3_2_A_X ),
    .C(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or3_2_C_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B2(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_B2_X ));
 sky130_fd_sc_hd__dfxtp_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[8] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net450),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net481),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.round_q[8] ),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.round_q[8] ),
    .A2(net451),
    .B1(net250),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_A ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .C(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o21a_2_A1_1_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_X ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_A_sky130_fd_sc_hd__o211a_2_X  (.A1(net451),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_A2 ),
    .B1(net401),
    .C1(net468),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_A ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1  (.A1(\m_blake2.m_hash256.round_q[8] ),
    .A2(net451),
    .A3(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X ),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1  (.A1(\m_blake2.m_hash256.round_q[8] ),
    .A2(net459),
    .A3(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(net444),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1 ),
    .B(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_C ),
    .D(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_X ));
 sky130_fd_sc_hd__o41a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__o41a_2_X  (.A1(net455),
    .A2(net459),
    .A3(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .A4(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_D_C ));
 sky130_fd_sc_hd__and3b_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__and3b_2_X  (.A_N(net468),
    .B(net469),
    .C(net474),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_X ),
    .C(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_C ),
    .D(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o211a_2_A2_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_C_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_C ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1 ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X ),
    .C(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_C ),
    .D(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_C_sky130_fd_sc_hd__o31a_2_X  (.A1(net458),
    .A2(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or2_2_B_X ),
    .A3(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(net444),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_C ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1  (.A1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o31a_2_B1_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.round_q[8] ),
    .B(net450),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B  (.A(net449),
    .B(\m_blake2.m_hash256.round_q[8] ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__or3_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.round_q[8] ),
    .B(net452),
    .C(net454),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1  (.A(\m_blake2.m_hash256.round_q[8] ),
    .B(net459),
    .C(net461),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o31a_2_A3  (.A1(net453),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .A3(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o31a_2_A3_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A  (.A(\m_blake2.m_hash256.round_q[8] ),
    .B(net450),
    .C(net457),
    .D(net462),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(net456),
    .A2(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(net444),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3  (.A1(net451),
    .A2(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A2_B1_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A3(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_1_X_sky130_fd_sc_hd__or4_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_2  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_2_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .B(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ));
 sky130_fd_sc_hd__nand2b_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B  (.A_N(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_1  (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__o31a_2_B1_X ),
    .B(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A_X ),
    .Y(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.round_q[9] ));
 sky130_fd_sc_hd__o211a_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_blake2.m_hash256.round_q[8] ),
    .A2(net152),
    .B1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net1710),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(net449),
    .B(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1  (.A1(net449),
    .A2(net455),
    .A3(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(net444),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1  (.A1(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_A2 ),
    .B1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X ),
    .C1(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__o211a_2_C1_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_X ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_A2_sky130_fd_sc_hd__or4_2_X  (.A(net455),
    .B(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ),
    .C(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .D(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__a211o_2_B1_A2 ));
 sky130_fd_sc_hd__or2_4 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A  (.A(net449),
    .B(net454),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A  (.A(\m_blake2.m_hash256.round_q[9] ),
    .B(net458),
    .C(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1  (.A(net449),
    .B(net450),
    .C(net453),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(net455),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_1_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2  (.A(net449),
    .B(net455),
    .C(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C_sky130_fd_sc_hd__or2_2_X  (.A(net457),
    .B(net459),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_C ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X_sky130_fd_sc_hd__o21a_2_A2  (.A1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X ),
    .B1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_2_X_sky130_fd_sc_hd__o21a_2_A2_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3  (.A(net449),
    .B(net457),
    .C(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X_sky130_fd_sc_hd__o31a_2_A3  (.A1(net453),
    .A2(net455),
    .A3(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X ),
    .B1(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_3_X_sky130_fd_sc_hd__o31a_2_A3_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_A2 ),
    .B1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X ),
    .B2(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o41a_2_A2_B1 ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_A2_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or3_2_A_X_sky130_fd_sc_hd__a22o_2_B1_A2 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A  (.A(net449),
    .B(net454),
    .C(net460),
    .D(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or3_2_A_1_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o31a_2_A1_B1 ),
    .A2(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X ),
    .B1(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_B1 ),
    .B2(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_B1_sky130_fd_sc_hd__or3_2_X  (.A(net407),
    .B(net458),
    .C(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .X(\m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_B1 ));
 sky130_fd_sc_hd__a21oi_4 \m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1  (.A1(net446),
    .A2(net478),
    .B1(net507),
    .Y(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(net852),
    .Q(\m_blake2.m_hash256.shift_hash_q ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net446),
    .A2(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A_Y ),
    .B1(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1 ),
    .Y(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(net446),
    .A2(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A_Y ),
    .B1(\m_blake2.m_hash256.fsm_q[5] ),
    .Y(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_io.cmd[5] ),
    .A2(\m_io.cmd[4] ),
    .B1(\m_blake2.m_hash256.slow_output_q ),
    .Y(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(net821),
    .Q(\m_blake2.m_hash256.slow_output_q ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(net820),
    .B(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__a21oi_2_B1_Y ),
    .Y(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A  (.A(net851),
    .Y(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[0][0] ),
    .A2(net402),
    .B1(\m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .C1(\m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .X(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .A2(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ),
    .B1(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .X(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1137),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][0] ),
    .B(\m_blake2.m_hash256.v_q[8][0] ),
    .X(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A2(\hash[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21oi_2_B1_Y ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C  (.A(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B(\hash[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .C(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][10] ),
    .A1(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ),
    .S(net363),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net401),
    .A2(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__o22a_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[11]_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__a21oi_2_Y_A1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net102),
    .B2(\m_blake2.m_hash256.m_matrix[0][10] ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][10] ),
    .A2(net146),
    .B1(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net107),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][10] ),
    .A2(net87),
    .B1(net111),
    .B2(\m_blake2.m_hash256.m_matrix[7][10] ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][10] ),
    .A2(net143),
    .B1(net99),
    .B2(\m_blake2.m_hash256.m_matrix[6][10] ),
    .C1(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][10] ),
    .A2(net127),
    .B1(net115),
    .B2(\m_blake2.m_hash256.m_matrix[5][10] ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][10] ),
    .A2(net91),
    .B1(net119),
    .B2(\m_blake2.m_hash256.m_matrix[13][10] ),
    .C1(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][10] ),
    .A2(net138),
    .B1(net95),
    .B2(\m_blake2.m_hash256.m_matrix[12][10] ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][10] ),
    .A2(net131),
    .B1(net151),
    .B2(\m_blake2.m_hash256.m_matrix[11][10] ),
    .C1(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][10] ),
    .A2(net135),
    .B1(net123),
    .B2(\m_blake2.m_hash256.m_matrix[15][10] ),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1010),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][10] ),
    .B(\m_blake2.m_hash256.v_q[8][10] ),
    .Y(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1513),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][11] ),
    .B(\m_blake2.m_hash256.v_q[8][11] ),
    .Y(\m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2  (.A1(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .A2(\m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1_N(net530),
    .X(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_B2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .B(\m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__o22a_2_A2_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][12] ),
    .A1(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .S(net372),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .A2(\m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net403),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__o22a_2 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][12] ),
    .A2(net100),
    .B1(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][12] ),
    .A2(net96),
    .B1(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net104),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][12] ),
    .A2(net108),
    .B1(net128),
    .B2(\m_blake2.m_hash256.m_matrix[8][12] ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][12] ),
    .A2(net116),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][12] ),
    .C1(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][12] ),
    .A2(net124),
    .B1(net112),
    .B2(\m_blake2.m_hash256.m_matrix[5][12] ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][12] ),
    .A2(net132),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][12] ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][12] ),
    .A2(net84),
    .B1(net88),
    .B2(\m_blake2.m_hash256.m_matrix[14][12] ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][12] ),
    .A2(net140),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][12] ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][12] ),
    .A2(net136),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][12] ),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1090),
    .S(net410),
    .X(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][12] ),
    .B(\m_blake2.m_hash256.v_q[8][12] ),
    .Y(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2  (.A1(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .A2(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1_N(net511),
    .X(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_B2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .B(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__o22a_2_A2_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1467),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][13] ),
    .B(\m_blake2.m_hash256.v_q[8][13] ),
    .Y(\m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B(\m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][14] ),
    .A1(\m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net386),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22oi_4 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2  (.A1(net404),
    .A2(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B2(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .Y(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ));
 sky130_fd_sc_hd__nand2b_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__nand2b_2_A_N  (.A_N(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ),
    .B(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A ),
    .Y(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and3_2_B_A ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net101),
    .B2(\m_blake2.m_hash256.m_matrix[0][14] ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][14] ),
    .A2(net129),
    .B1(net97),
    .B2(\m_blake2.m_hash256.m_matrix[6][14] ),
    .C1(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][14] ),
    .A2(net137),
    .B1(net117),
    .B2(\m_blake2.m_hash256.m_matrix[13][14] ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][14] ),
    .A2(net85),
    .B1(net113),
    .B2(\m_blake2.m_hash256.m_matrix[5][14] ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][14] ),
    .A2(net89),
    .B1(net145),
    .B2(\m_blake2.m_hash256.m_matrix[10][14] ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][14] ),
    .A2(net109),
    .B1(net121),
    .B2(\m_blake2.m_hash256.m_matrix[15][14] ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][14] ),
    .A2(net125),
    .B1(net105),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][14] ),
    .A2(net141),
    .B1(net93),
    .B2(\m_blake2.m_hash256.m_matrix[12][14] ),
    .C1(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][14] ),
    .A2(net133),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][14] ),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1111),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][14] ),
    .B(\m_blake2.m_hash256.v_q[8][14] ),
    .Y(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][15] ),
    .A1(\m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net389),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_2 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net404),
    .A2(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B2(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .X(\m_blake2.m_hash256.m_g.a0[16]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__nor3_2_Y_A ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][15] ),
    .A2(net101),
    .B1(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][15] ),
    .A2(net125),
    .B1(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net105),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][15] ),
    .A2(net145),
    .B1(net97),
    .B2(\m_blake2.m_hash256.m_matrix[6][15] ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][15] ),
    .A2(net117),
    .B1(net93),
    .B2(\m_blake2.m_hash256.m_matrix[12][15] ),
    .C1(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][15] ),
    .A2(net129),
    .B1(net133),
    .B2(\m_blake2.m_hash256.m_matrix[3][15] ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][15] ),
    .A2(net137),
    .B1(net121),
    .B2(\m_blake2.m_hash256.m_matrix[15][15] ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][15] ),
    .A2(net85),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][15] ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][15] ),
    .A2(net109),
    .B1(net141),
    .B2(\m_blake2.m_hash256.m_matrix[1][15] ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][15] ),
    .A2(net89),
    .B1(net113),
    .B2(\m_blake2.m_hash256.m_matrix[5][15] ),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .Y(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1040),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][15] ),
    .B(\m_blake2.m_hash256.v_q[8][15] ),
    .Y(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][16] ),
    .A1(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net362),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .A2(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_A2 ),
    .B1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net402),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A ),
    .A2(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B ),
    .B1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A ),
    .B(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B ),
    .C(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][16] ),
    .B(net103),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A ));
 sky130_fd_sc_hd__or3_4 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X  (.A(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B ),
    .C(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][16] ),
    .A2(net134),
    .B1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][16] ),
    .A2(net118),
    .B1(net94),
    .B2(\m_blake2.m_hash256.m_matrix[12][16] ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][16] ),
    .A2(net86),
    .B1(net98),
    .B2(\m_blake2.m_hash256.m_matrix[6][16] ),
    .C1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][16] ),
    .A2(net110),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][16] ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][16] ),
    .A2(net130),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][16] ),
    .C1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][16] ),
    .A2(net138),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][16] ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][16] ),
    .A2(net114),
    .B1(net146),
    .B2(\m_blake2.m_hash256.m_matrix[10][16] ),
    .C1(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][16] ),
    .A2(net126),
    .B1(net90),
    .B2(\m_blake2.m_hash256.m_matrix[14][16] ),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net980),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][16] ),
    .B(\m_blake2.m_hash256.v_q[8][16] ),
    .Y(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][17] ),
    .A1(\m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net362),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ),
    .A2(\m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net402),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net100),
    .B2(\m_blake2.m_hash256.m_matrix[0][17] ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][17] ),
    .A2(net114),
    .B1(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][17] ),
    .A2(net90),
    .B1(net146),
    .B2(\m_blake2.m_hash256.m_matrix[10][17] ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][17] ),
    .A2(net118),
    .B1(net98),
    .B2(\m_blake2.m_hash256.m_matrix[6][17] ),
    .C1(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][17] ),
    .A2(net94),
    .B1(net150),
    .B2(\m_blake2.m_hash256.m_matrix[11][17] ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][17] ),
    .A2(net138),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][17] ),
    .C1(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][17] ),
    .A2(net126),
    .B1(net86),
    .B2(\m_blake2.m_hash256.m_matrix[4][17] ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][17] ),
    .A2(net110),
    .B1(net130),
    .B2(\m_blake2.m_hash256.m_matrix[8][17] ),
    .C1(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][17] ),
    .A2(net134),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][17] ),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net914),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][17] ),
    .B(\m_blake2.m_hash256.v_q[8][17] ),
    .Y(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][18] ),
    .A1(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net363),
    .X(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_Y ),
    .A2(\m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net402),
    .X(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1  (.A1(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_A ),
    .A2(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B ),
    .B1(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net970),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][18] ),
    .B(\m_blake2.m_hash256.v_q[8][18] ),
    .Y(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[18]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][19] ),
    .A1(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net390),
    .X(\m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_2 \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net405),
    .A2(\m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B2(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .A1(net1058),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][19] ),
    .B(\m_blake2.m_hash256.v_q[8][19] ),
    .Y(\m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net998),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][1] ),
    .A1(\hash[1]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .S(net363),
    .X(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .A2(\m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net402),
    .X(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][1] ),
    .B(\m_blake2.m_hash256.v_q[8][1] ),
    .Y(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\hash[1]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .B(\m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[9]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][20] ),
    .A1(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net372),
    .X(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_X ),
    .A2(\m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net403),
    .X(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net960),
    .S(net410),
    .X(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][20] ),
    .B(\m_blake2.m_hash256.v_q[8][20] ),
    .Y(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][21] ),
    .A1(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net378),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(\m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__a211oi_2_A1_Y ),
    .A2_N(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ),
    .B1(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net406),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[22]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net100),
    .B2(\m_blake2.m_hash256.m_matrix[0][21] ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][21] ),
    .A2(net108),
    .B1(net128),
    .B2(\m_blake2.m_hash256.m_matrix[8][21] ),
    .C1(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][21] ),
    .A2(net88),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][21] ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][21] ),
    .A2(net132),
    .B1(net136),
    .B2(\m_blake2.m_hash256.m_matrix[2][21] ),
    .C1(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][21] ),
    .A2(net84),
    .B1(net140),
    .B2(\m_blake2.m_hash256.m_matrix[1][21] ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][21] ),
    .A2(net112),
    .B1(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net104),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][21] ),
    .A2(net92),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][21] ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][21] ),
    .A2(net116),
    .B1(net96),
    .B2(\m_blake2.m_hash256.m_matrix[6][21] ),
    .C1(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][21] ),
    .A2(net124),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][21] ),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1052),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][21] ),
    .B(\m_blake2.m_hash256.v_q[8][21] ),
    .Y(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][22] ),
    .A1(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net386),
    .X(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_2 \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_X ),
    .A2(\m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net404),
    .X(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ),
    .C(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net993),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][22] ),
    .B(\m_blake2.m_hash256.v_q[8][22] ),
    .Y(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][23] ),
    .A1(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net389),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_2 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .A2(\m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net404),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o32a_2 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net101),
    .B2(\m_blake2.m_hash256.m_matrix[0][23] ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][23] ),
    .A2(net125),
    .B1(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net105),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][23] ),
    .A2(net129),
    .B1(net137),
    .B2(\m_blake2.m_hash256.m_matrix[2][23] ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][23] ),
    .A2(net85),
    .B1(net121),
    .B2(\m_blake2.m_hash256.m_matrix[15][23] ),
    .C1(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][23] ),
    .A2(net89),
    .B1(net93),
    .B2(\m_blake2.m_hash256.m_matrix[12][23] ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[10][23] ),
    .A2(net145),
    .B1(net97),
    .B2(\m_blake2.m_hash256.m_matrix[6][23] ),
    .C1(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][23] ),
    .A2(net141),
    .B1(net117),
    .B2(\m_blake2.m_hash256.m_matrix[13][23] ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][23] ),
    .A2(net113),
    .B1(net133),
    .B2(\m_blake2.m_hash256.m_matrix[3][23] ),
    .C1(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][23] ),
    .A2(net109),
    .B1(net149),
    .B2(\m_blake2.m_hash256.m_matrix[11][23] ),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1093),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][23] ),
    .B(\m_blake2.m_hash256.v_q[8][23] ),
    .Y(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[23]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][24] ),
    .A1(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net372),
    .X(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22oi_4 \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2  (.A1(net403),
    .A2(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B2(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .Y(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .A1(net1127),
    .S(net410),
    .X(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][24] ),
    .B(\m_blake2.m_hash256.v_q[8][24] ),
    .Y(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][25] ),
    .A1(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net366),
    .X(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net402),
    .A2(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B2(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .X(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N ),
    .B(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .Y(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1085),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][25] ),
    .B(\m_blake2.m_hash256.v_q[8][25] ),
    .Y(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][26] ),
    .A1(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net367),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B  (.A(net401),
    .B(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1  (.A1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ),
    .A2(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2 ),
    .B1(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .C1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_X ));
 sky130_fd_sc_hd__or2_2 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.m_matrix[0][26] ),
    .B(net102),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ));
 sky130_fd_sc_hd__or3_2 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X  (.A(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B ),
    .C(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][26] ),
    .A2(net87),
    .B1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net106),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][26] ),
    .A2(net115),
    .B1(net147),
    .B2(\m_blake2.m_hash256.m_matrix[10][26] ),
    .C1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][26] ),
    .A2(net110),
    .B1(net122),
    .B2(\m_blake2.m_hash256.m_matrix[15][26] ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][26] ),
    .A2(net135),
    .B1(net119),
    .B2(\m_blake2.m_hash256.m_matrix[13][26] ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][26] ),
    .A2(net127),
    .B1(net98),
    .B2(\m_blake2.m_hash256.m_matrix[6][26] ),
    .C1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][26] ),
    .A2(net90),
    .B1(net130),
    .B2(\m_blake2.m_hash256.m_matrix[8][26] ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[12][26] ),
    .A2(net95),
    .B1(net151),
    .B2(\m_blake2.m_hash256.m_matrix[11][26] ),
    .C1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][26] ),
    .A2(net138),
    .B1(net142),
    .B2(\m_blake2.m_hash256.m_matrix[1][26] ),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__o211ai_4 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__o211ai_2_A2  (.A1(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .A2(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X ),
    .B1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A1 ),
    .C1(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2 ),
    .Y(\m_blake2.m_hash256.m_g.a0[27]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and3_2_X_A ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net973),
    .S(net410),
    .X(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][26] ),
    .B(\m_blake2.m_hash256.v_q[8][26] ),
    .Y(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][27] ),
    .A1(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net390),
    .X(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_2 \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2  (.A1_N(\m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__a211oi_2_A1_Y ),
    .A2_N(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ),
    .B1(net405),
    .B2(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .X(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2 ),
    .B(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X ),
    .Y(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net967),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][27] ),
    .B(\m_blake2.m_hash256.v_q[8][27] ),
    .Y(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[27]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][28] ),
    .A1(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net378),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .A2(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_A2 ),
    .B1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net406),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B  (.A(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o22a_4 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X  (.A1(\m_blake2.m_hash256.m_matrix[0][28] ),
    .A2(net100),
    .B1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ),
    .B2(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][28] ),
    .A2(net136),
    .B1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net104),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][28] ),
    .A2(net108),
    .B1(net112),
    .B2(\m_blake2.m_hash256.m_matrix[5][28] ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][28] ),
    .A2(net96),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][28] ),
    .C1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][28] ),
    .A2(net132),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][28] ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__or4_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X  (.A(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ),
    .C(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ),
    .D(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][28] ),
    .A2(net84),
    .B1(net116),
    .B2(\m_blake2.m_hash256.m_matrix[13][28] ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][28] ),
    .A2(net124),
    .B1(net128),
    .B2(\m_blake2.m_hash256.m_matrix[8][28] ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][28] ),
    .A2(net140),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][28] ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[14][28] ),
    .A2(net88),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][28] ),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B  (.A(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net949),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][28] ),
    .B(\m_blake2.m_hash256.v_q[8][28] ),
    .Y(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][29] ),
    .A1(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net385),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__o2bb2a_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N  (.A1_N(net404),
    .A2_N(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__a211oi_2_A1_Y ),
    .B2(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_X ),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ),
    .Y(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X ),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_A ));
 sky130_fd_sc_hd__a32o_4 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X  (.A1(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1 ),
    .A2(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2 ),
    .A3(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3 ),
    .B1(net104),
    .B2(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_B2 ),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__a221oi_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y  (.A1(\m_blake2.m_hash256.m_matrix[4][29] ),
    .A2(net84),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][29] ),
    .C1(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1 ),
    .Y(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[2][29] ),
    .A2(net136),
    .B1(net140),
    .B2(\m_blake2.m_hash256.m_matrix[1][29] ),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1 ));
 sky130_fd_sc_hd__a2111oi_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y  (.A1(\m_blake2.m_hash256.m_matrix[11][29] ),
    .A2(net148),
    .B1(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1 ),
    .D1(net104),
    .Y(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[3][29] ),
    .A2(net132),
    .B1(net96),
    .B2(\m_blake2.m_hash256.m_matrix[6][29] ),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][29] ),
    .A2(net108),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][29] ),
    .C1(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][29] ),
    .A2(net128),
    .B1(net112),
    .B2(\m_blake2.m_hash256.m_matrix[5][29] ),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221oi_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y  (.A1(\m_blake2.m_hash256.m_matrix[14][29] ),
    .A2(net88),
    .B1(net116),
    .B2(\m_blake2.m_hash256.m_matrix[13][29] ),
    .C1(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1 ),
    .Y(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][29] ),
    .A2(net124),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][29] ),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1 ));
 sky130_fd_sc_hd__inv_2 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_B2_sky130_fd_sc_hd__inv_2_Y  (.A(\m_blake2.m_hash256.m_matrix[0][29] ),
    .Y(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_B2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ),
    .A1(net1272),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][29] ),
    .B(\m_blake2.m_hash256.v_q[8][29] ),
    .Y(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1290),
    .S(net410),
    .X(\m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][2] ),
    .B(\m_blake2.m_hash256.v_q[8][2] ),
    .Y(\m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\hash[2]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .B(\m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[10]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][30] ),
    .A1(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net389),
    .X(\m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net404),
    .A2(\m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B2(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1048),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][30] ),
    .B(\m_blake2.m_hash256.v_q[8][30] ),
    .Y(\m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[30]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][31] ),
    .A1(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net390),
    .X(\m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(\m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__a211oi_2_A1_Y ),
    .A2_N(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_Y ),
    .B1(\m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net404),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net990),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][31] ),
    .B(\m_blake2.m_hash256.v_q[8][31] ),
    .Y(\m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[31]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net984),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][3] ),
    .A1(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .S(net392),
    .X(\m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_2 \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .A2(\m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net405),
    .X(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_A2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][3] ),
    .B(\m_blake2.m_hash256.v_q[8][3] ),
    .Y(\m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2  (.A1(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A2(\m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1_N(net531),
    .X(\m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2_B2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B(\m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1405),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][4] ),
    .B(\m_blake2.m_hash256.v_q[8][4] ),
    .Y(\m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2  (.A1(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .A2(\m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1_N(net510),
    .X(\m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2_B2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B(\m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net950),
    .S(net412),
    .X(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][5] ),
    .A1(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .S(net379),
    .X(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1  (.A1(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .A2(\m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net404),
    .X(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][5] ),
    .B(\m_blake2.m_hash256.v_q[8][5] ),
    .Y(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2  (.A1(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .A2(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1_N(net517),
    .X(\m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2_B2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .B(\m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net974),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][6] ),
    .A1(\hash[6]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net386),
    .X(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2  (.A1(net404),
    .A2(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .B2(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_X ),
    .X(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][6] ),
    .B(\m_blake2.m_hash256.v_q[8][6] ),
    .Y(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\hash[6]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net991),
    .S(net411),
    .X(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][7] ),
    .A1(\hash[7]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net391),
    .X(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a21o_2 \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net404),
    .A2(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][7] ),
    .B(\m_blake2.m_hash256.v_q[8][7] ),
    .Y(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\hash[7]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .A1(net1254),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[0][8] ),
    .A1(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .S(net366),
    .X(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_Y ),
    .A2_N(\m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__a211oi_2_A1_Y ),
    .B1(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net402),
    .X(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__and2b_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ),
    .B(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][8] ),
    .B(\m_blake2.m_hash256.v_q[8][8] ),
    .Y(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__a21bo_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2  (.A1(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .A2(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B1_N(net501),
    .X(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__o22a_2_A2_B2 ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B  (.A(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .B(\m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[16]_sky130_fd_sc_hd__o22a_2_A2_B1 ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[0][9] ),
    .A2(net402),
    .B1(\m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .C1(\m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .Y(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1  (.A1(net363),
    .A2(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .A3(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y ),
    .X(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1_X ));
 sky130_fd_sc_hd__a211oi_2 \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__a211oi_2_C1  (.A1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1 ),
    .A2(net105),
    .B1(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ),
    .C1(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_Y_sky130_fd_sc_hd__a31o_2_B1_X ),
    .Y(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor3_2_B_A ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[0][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1414),
    .S(net409),
    .X(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[0][9] ),
    .B(\m_blake2.m_hash256.v_q[8][9] ),
    .Y(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B(\m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[17]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][0] ),
    .A2(net169),
    .B1(net171),
    .B2(\m_blake2.m_hash256.v_q[11][0] ),
    .X(\m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1712),
    .A1(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][10] ),
    .A2(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ),
    .B1(\m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net171),
    .C1(\m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.g_c_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1777),
    .A1(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1000),
    .A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[10][11] ),
    .B(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ),
    .Y(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__and3_4 \m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X  (.A(net408),
    .B(net355),
    .C(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1211),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net234),
    .X(\m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][12] ),
    .A2(net372),
    .B1(net169),
    .X(\m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1377),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][13] ),
    .A2(net378),
    .B1(net169),
    .X(\m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[10][14] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][14] ),
    .A2(net379),
    .B1(net407),
    .X(\m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1631),
    .A1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][15] ),
    .A2(net386),
    .B1(net170),
    .X(\m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][16] ),
    .A2(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ),
    .B1(\m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net171),
    .C1(\m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.g_c_buf[16]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1064),
    .A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1745),
    .A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][17] ),
    .A2(net365),
    .B1(net169),
    .X(\m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_D1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[10][18] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][18] ),
    .A2(net364),
    .B1(net169),
    .X(\m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_D1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1665),
    .A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][19] ),
    .A2(net388),
    .B1(net408),
    .X(\m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net916),
    .A1(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[10][1] ),
    .B(net364),
    .X(\m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[10][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1105),
    .A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net234),
    .X(\m_blake2.m_hash256.v_q[10][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net876),
    .A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[10][21] ),
    .B(net379),
    .X(\m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1527),
    .A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][22] ),
    .A2(net387),
    .B1(net170),
    .X(\m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[10][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1772),
    .A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[10][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1300),
    .A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net234),
    .X(\m_blake2.m_hash256.v_q[10][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][25] ),
    .A2(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ),
    .B1(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_X ),
    .B2(net249),
    .X(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1324),
    .A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1902),
    .A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][26] ),
    .A2(net367),
    .B1(net169),
    .X(\m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1874),
    .A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[10][27] ),
    .B(net391),
    .X(\m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net958),
    .A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[10][28] ),
    .B(net378),
    .X(\m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1083),
    .A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][29] ),
    .A2(net386),
    .B1(net170),
    .X(\m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][2] ),
    .A2(net169),
    .B1(net171),
    .B2(\m_blake2.m_hash256.v_q[11][2] ),
    .X(\m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1263),
    .A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net234),
    .X(\m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B  (.A(net408),
    .B(\m_blake2.m_hash256.v_q[10][30] ),
    .C(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B  (.A(net477),
    .B(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .Y(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1  (.A(net407),
    .B(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .Y(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1_Y ));
 sky130_fd_sc_hd__xor2_4 \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__xor2_2_X  (.A(net466),
    .B(net471),
    .X(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1233),
    .A1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.v_q[10][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[10][31] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[10][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1820),
    .A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1023),
    .A1(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[10][4] ),
    .B(net378),
    .X(\m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1351),
    .A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__o31a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][5] ),
    .A2(net385),
    .A3(net249),
    .B1(net408),
    .X(\m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1306),
    .A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net235),
    .X(\m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][6] ),
    .A2(net387),
    .B1(net170),
    .X(\m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][7] ),
    .A2(net170),
    .B1(net172),
    .B2(\m_blake2.m_hash256.v_q[11][7] ),
    .X(\m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[10][7] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net236),
    .X(\m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1411),
    .A1(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][8] ),
    .A2(net366),
    .B1(net169),
    .X(\m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[10][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[10][9] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net233),
    .X(\m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[10][9] ),
    .A2(net362),
    .B1(net407),
    .X(\m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[11][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][0]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1584),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .A1(net1543),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][10] ),
    .B(net364),
    .X(\m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[11][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1330),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .A1(net1395),
    .S(net218),
    .X(\m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][12] ),
    .B(net372),
    .X(\m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1460),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__o22a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][13] ),
    .A2(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ),
    .B1(net173),
    .B2(net254),
    .X(\m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1656),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][14] ),
    .A2(net379),
    .B1(net172),
    .X(\m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(\m_blake2.m_hash256.v_q[11][15] ),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__o22a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][15] ),
    .A2(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ),
    .B1(net172),
    .B2(net253),
    .X(\m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .A1(net1801),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][16] ),
    .B(net362),
    .X(\m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1551),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][17] ),
    .A2(net362),
    .B1(net171),
    .X(\m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .A1(net1900),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][18] ),
    .A2(net364),
    .B1(net171),
    .X(\m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1867),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][19] ),
    .A2(net388),
    .B1(net173),
    .X(\m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1562),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][1] ),
    .A2(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ),
    .B1(net171),
    .B2(net254),
    .X(\m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__or2_4 \m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2_sky130_fd_sc_hd__or2_2_X  (.A(net362),
    .B(net254),
    .X(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[11][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .A1(net1065),
    .S(net218),
    .X(\m_blake2.m_hash256.v_q[11][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[11][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1681),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1614),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][22] ),
    .A2(net387),
    .B1(net172),
    .X(\m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][23] ),
    .A2(net172),
    .B1(\m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__a22o_2_B1_X ),
    .C1(net253),
    .X(\m_blake2.m_hash256.g_c_buf[23]_sky130_fd_sc_hd__o311a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(\m_blake2.m_hash256.v_q[11][23] ),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .A1(net1082),
    .S(net218),
    .X(\m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][24] ),
    .B(net372),
    .X(\m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[11][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1735),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1697),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][26] ),
    .B(net367),
    .X(\m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][27] ),
    .A2(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net408),
    .X(\m_blake2.m_hash256.g_c_buf[27]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(\m_blake2.m_hash256.v_q[11][27] ),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[11][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1112),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1275),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__o22a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][29] ),
    .A2(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ),
    .B1(net172),
    .B2(net253),
    .X(\m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[11][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][2]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1849),
    .S(net218),
    .X(\m_blake2.m_hash256.v_q[11][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[11][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1626),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1817),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][31] ),
    .B(net388),
    .X(\m_blake2.m_hash256.v_q[11][31]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1430),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][3] ),
    .B(net393),
    .X(\m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1507),
    .S(net220),
    .X(\m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][4] ),
    .A2(net378),
    .B1(net173),
    .X(\m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1742),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][5] ),
    .A2(net385),
    .B1(net172),
    .X(\m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[11][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][6]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1762),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[11][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][7]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(\m_blake2.m_hash256.v_q[11][7] ),
    .S(net219),
    .X(\m_blake2.m_hash256.v_q[11][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .A1(net1252),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[11][8] ),
    .B(net366),
    .X(\m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[11][9] ),
    .A2(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ),
    .B1(\m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net250),
    .C1(\m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.g_c_buf[9]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[11][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(\m_blake2.m_hash256.v_q[11][9] ),
    .S(net217),
    .X(\m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[12][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][0]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1542),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][10] ),
    .A2(net344),
    .B1(net259),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[4] ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1486),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][11] ),
    .A2(net350),
    .B1(net260),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[5] ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .A1(net1161),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1598),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][12] ),
    .B(net352),
    .Y(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[12][13] ),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[12][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1783),
    .S(net228),
    .X(\m_blake2.m_hash256.v_q[12][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][14]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][14] ),
    .B(net353),
    .Y(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[12][15] ),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1718),
    .S(net226),
    .X(\m_blake2.m_hash256.v_q[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1861),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][17] ),
    .B(net343),
    .Y(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1271),
    .S(net226),
    .X(\m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][18] ),
    .B(net347),
    .Y(\m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[12][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1349),
    .S(net226),
    .X(\m_blake2.m_hash256.v_q[12][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][19]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][19] ),
    .B(net347),
    .Y(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[12][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][1]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1829),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.v_q[12][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1600),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][21] ),
    .A2(net358),
    .B1(net262),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[15] ),
    .C1(net269),
    .X(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[12][21] ),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][22]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][22] ),
    .A2(net351),
    .B1(net263),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[16] ),
    .C1(net269),
    .X(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[12][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1780),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][23] ),
    .A2(net357),
    .B1(net261),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[17] ),
    .C1(net269),
    .X(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(\m_blake2.m_hash256.v_q[12][23] ),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1493),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][24] ),
    .B(net349),
    .Y(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[12][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1798),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1321),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][27] ),
    .A2(net349),
    .B1(net260),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[21] ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1373),
    .S(net226),
    .X(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1541),
    .S(net228),
    .X(\m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][28] ),
    .B(net353),
    .Y(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][29] ),
    .A2(net358),
    .B1(net262),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[23] ),
    .C1(net269),
    .X(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1869),
    .S(net228),
    .X(\m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[12][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][2]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1632),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[12][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1845),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][30]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][30] ),
    .B(net357),
    .Y(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1879),
    .S(net228),
    .X(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1683),
    .S(net228),
    .X(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net983),
    .S(net228),
    .X(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1466),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1770),
    .S(net228),
    .X(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][6] ),
    .B(net351),
    .Y(\m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[12][7] ),
    .S(net227),
    .X(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[12][8] ),
    .A2(net347),
    .B1(net260),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[2] ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1763),
    .S(net226),
    .X(\m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[12][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1653),
    .S(net225),
    .X(\m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[12][9] ),
    .B(net343),
    .Y(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][0]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][0] ),
    .A2(net347),
    .B1(net259),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[26] ),
    .C1(\m_io.m_config.ll_q[32]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[13][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][0]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1412),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][10] ),
    .A2(net347),
    .B1(net260),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[36] ),
    .C1(\m_io.m_config.ll_q[42]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1443),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .A1(net1658),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.v_q[13][11] ),
    .B(net377),
    .Y(\m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][12] ),
    .A2(net357),
    .B1(net262),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[38] ),
    .C1(\m_io.m_config.ll_q[44]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1897),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[13][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[13][13] ),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__a2bb2o_2_A1_N  (.A1_N(\m_blake2.m_hash256.v_q[13][14] ),
    .A2_N(net380),
    .B1(net264),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[40] ),
    .X(\m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1182),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][15]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][15] ),
    .A2(net357),
    .B1(net261),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[41] ),
    .C1(\m_io.m_config.ll_q[47]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[13][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[13][15] ),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.v_q[13][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1550),
    .S(net208),
    .X(\m_blake2.m_hash256.v_q[13][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][17] ),
    .A2(net343),
    .B1(net259),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[43] ),
    .C1(\m_io.m_config.ll_q[49]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1842),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[13][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1372),
    .S(net208),
    .X(\m_blake2.m_hash256.v_q[13][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ba_1 \m_blake2.m_hash256.v_q[13][18]_sky130_fd_sc_hd__o21ba_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][18] ),
    .A2(net373),
    .B1_N(\m_io.m_config.ll_q[50]_sky130_fd_sc_hd__a22o_2_B2_X ),
    .X(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][19] ),
    .A2(net348),
    .B1(net260),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[45] ),
    .C1(\m_io.m_config.ll_q[51]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1622),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][1] ),
    .A2(net343),
    .B1(net259),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[27] ),
    .C1(\m_io.m_config.ll_q[33]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1876),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][20]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][20] ),
    .A2(net358),
    .B1(net261),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[46] ),
    .C1(\m_io.m_config.ll_q[52]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[13][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1613),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][21]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][21] ),
    .A2(net358),
    .B1(net262),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[47] ),
    .C1(\m_io.m_config.ll_q[53]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[13][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[13][21] ),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][22]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][22] ),
    .A2(net351),
    .B1(net263),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[48] ),
    .C1(\m_io.m_config.ll_q[54]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[13][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1247),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][23]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][23] ),
    .A2(net358),
    .B1(net261),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[49] ),
    .C1(\m_io.m_config.ll_q[55]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[13][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(\m_blake2.m_hash256.v_q[13][23] ),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__a2bb2o_2_A1_N  (.A1_N(\m_blake2.m_hash256.v_q[13][24] ),
    .A2_N(net380),
    .B1(net264),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[50] ),
    .X(\m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net920),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1816),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.v_q[13][25] ),
    .B(net368),
    .Y(\m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][26] ),
    .A2(net348),
    .B1(net260),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[52] ),
    .C1(\m_io.m_config.ll_q[58]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1577),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1659),
    .S(net208),
    .X(\m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_blake2.m_hash256.v_q[13][27] ),
    .B(net375),
    .Y(\m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__a2bb2o_2_A1_N  (.A1_N(\m_blake2.m_hash256.v_q[13][28] ),
    .A2_N(net382),
    .B1(net264),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[54] ),
    .X(\m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1026),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][29] ),
    .A2(net358),
    .B1(net262),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[55] ),
    .C1(\m_io.m_config.ll_q[61]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(\m_blake2.m_hash256.v_q[13][29] ),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[13][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][2]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1359),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][30]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][30] ),
    .A2(net357),
    .B1(net261),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[56] ),
    .C1(\m_io.m_config.ll_q[62]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[13][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1504),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[13][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1854),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.v_q[13][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][3]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1444),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][4]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][4] ),
    .A2(net352),
    .B1(net264),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[30] ),
    .C1(\m_io.m_config.ll_q[36]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.v_q[13][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][4]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1860),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][5]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][5] ),
    .A2(net358),
    .B1(net262),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[31] ),
    .C1(\m_io.m_config.ll_q[37]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[13][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][5]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[13][5] ),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][6] ),
    .A2(net351),
    .B1(net263),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[32] ),
    .C1(\m_io.m_config.ll_q[38]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__a221o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(net1567),
    .S(net207),
    .X(\m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[13][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][7]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .A1(\m_blake2.m_hash256.v_q[13][7] ),
    .S(net206),
    .X(\m_blake2.m_hash256.v_q[13][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][8] ),
    .A2(net349),
    .B1(net260),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[34] ),
    .C1(\m_io.m_config.ll_q[40]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1144),
    .S(net208),
    .X(\m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[13][9] ),
    .A2(net343),
    .B1(net259),
    .B2(\m_blake2.m_hash256.block_idx_plus_one_q[35] ),
    .C1(\m_io.m_config.ll_q[41]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[13][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1853),
    .S(net205),
    .X(\m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[14][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][0]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1307),
    .A1(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1366),
    .A1(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][10] ),
    .B(net369),
    .X(\m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.v_q[14][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1238),
    .A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .S(net212),
    .X(\m_blake2.m_hash256.v_q[14][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1007),
    .A1(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][12] ),
    .B(net394),
    .X(\m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[14][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[14][13] ),
    .A1(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][13]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][13] ),
    .B(net394),
    .X(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1029),
    .A1(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[14][14] ),
    .A2(net382),
    .B1(net186),
    .Y(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[14][15] ),
    .A1(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][15] ),
    .B(net393),
    .X(\m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[14][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net861),
    .A1(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][16]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][16] ),
    .B(net380),
    .X(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1678),
    .A1(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][17] ),
    .B(net369),
    .X(\m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[14][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1608),
    .A1(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net212),
    .X(\m_blake2.m_hash256.v_q[14][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1024),
    .A1(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][19] ),
    .B(net373),
    .X(\m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[14][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][1]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[14][1] ),
    .A1(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net910),
    .A1(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][20] ),
    .B(net395),
    .X(\m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[14][21] ),
    .A1(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][21] ),
    .B(net394),
    .X(\m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1022),
    .A1(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][22] ),
    .B(net383),
    .X(\m_blake2.m_hash256.v_q[14][22]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[14][23] ),
    .A1(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][23] ),
    .B(net393),
    .X(\m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1299),
    .A1(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[14][24] ),
    .A2(net380),
    .B1(net186),
    .Y(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[14][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1575),
    .A1(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1154),
    .A1(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][26] ),
    .B(net373),
    .X(\m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[14][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net943),
    .A1(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net212),
    .X(\m_blake2.m_hash256.v_q[14][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1458),
    .A1(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[14][28] ),
    .A2(net382),
    .B1(net186),
    .Y(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1749),
    .A1(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][29] ),
    .B(net394),
    .X(\m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[14][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][2]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1457),
    .A1(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1018),
    .A1(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][30] ),
    .B(net392),
    .X(\m_blake2.m_hash256.v_q[14][30]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[14][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1173),
    .A1(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][31]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][31] ),
    .B(net392),
    .X(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_blake2.m_hash256.v_q[14][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1596),
    .A1(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[14][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][4]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1092),
    .A1(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[14][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][5]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[14][5] ),
    .A1(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1352),
    .A1(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net211),
    .X(\m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][6] ),
    .B(net383),
    .X(\m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[14][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][7]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1727),
    .A1(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net210),
    .X(\m_blake2.m_hash256.v_q[14][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][7]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][7] ),
    .B(net393),
    .X(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1125),
    .A1(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][8] ),
    .B(net376),
    .X(\m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[14][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1785),
    .A1(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net209),
    .X(\m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[14][9] ),
    .B(net369),
    .X(\m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[15][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][0]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1011),
    .A1(\m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net858),
    .A1(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[15][10] ),
    .B(net369),
    .X(\m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1314),
    .A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .S(net297),
    .X(\m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][11] ),
    .A2(net377),
    .B1(net193),
    .Y(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][12] ),
    .A2(net276),
    .B1(\m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net186),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1169),
    .A1(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[15][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1733),
    .A1(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1320),
    .A1(\m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net299),
    .X(\m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][14] ),
    .A2(net382),
    .B1(net194),
    .Y(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1322),
    .A1(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[15][15] ),
    .B(net393),
    .X(\m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[15][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1207),
    .A1(\m_blake2.m_hash256.m_g.d_q[8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net297),
    .X(\m_blake2.m_hash256.v_q[15][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][17] ),
    .A2(net275),
    .B1(\m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net185),
    .C1(net270),
    .X(\m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1654),
    .A1(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[15][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1147),
    .A1(\m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net297),
    .X(\m_blake2.m_hash256.v_q[15][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][19] ),
    .A2(net275),
    .B1(net176),
    .B2(\m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__or2_2_A_X ),
    .C1(net271),
    .X(\m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1441),
    .A1(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[15][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][1]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1295),
    .A1(\m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][20] ),
    .A2(net276),
    .B1(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__or2_2_A_X ),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1435),
    .A1(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1509),
    .A1(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net299),
    .X(\m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[15][21] ),
    .B(net394),
    .X(\m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net898),
    .A1(\m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[15][22] ),
    .B(net383),
    .X(\m_blake2.m_hash256.v_q[15][22]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1388),
    .A1(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[15][23] ),
    .B(net392),
    .X(\m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1120),
    .A1(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net297),
    .X(\m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][24] ),
    .A2(net380),
    .B1(net193),
    .Y(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1213),
    .A1(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][25] ),
    .A2(net368),
    .B1(net193),
    .Y(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][26] ),
    .A2(net275),
    .B1(\m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net185),
    .C1(net271),
    .X(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1230),
    .A1(\m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[15][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1195),
    .A1(\m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net297),
    .X(\m_blake2.m_hash256.v_q[15][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[15][27]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][27] ),
    .A2(net375),
    .B1(net193),
    .Y(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1167),
    .A1(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net299),
    .X(\m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][28] ),
    .A2(net381),
    .B1(net194),
    .Y(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_C ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][29] ),
    .A2(net276),
    .B1(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ),
    .B2(\m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__or2_2_A_X ),
    .C1(net272),
    .X(\m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1809),
    .A1(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][2]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1218),
    .A1(\m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net824),
    .A1(\m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net299),
    .X(\m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[15][30] ),
    .B(net392),
    .X(\m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[15][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1442),
    .A1(\m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.v_q[15][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1451),
    .A1(\m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net299),
    .X(\m_blake2.m_hash256.v_q[15][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[15][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][4]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1448),
    .A1(\m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net299),
    .X(\m_blake2.m_hash256.v_q[15][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[15][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][5]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1690),
    .A1(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[15][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][6]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1170),
    .A1(\m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net299),
    .X(\m_blake2.m_hash256.v_q[15][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[15][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][7]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1669),
    .A1(\m_blake2.m_hash256.v_q[12][7]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net298),
    .X(\m_blake2.m_hash256.v_q[15][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net882),
    .A1(\m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[15][8] ),
    .B(net376),
    .X(\m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[15][9] ),
    .A2(net275),
    .B1(net176),
    .B2(\m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__or2_2_A_X ),
    .C1(net270),
    .X(\m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__nor2_4 \m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y  (.A(net259),
    .B(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[15][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1825),
    .A1(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net296),
    .X(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][0] ),
    .A2(net290),
    .B1(net278),
    .B2(\m_blake2.m_hash256.v_q[2][0] ),
    .X(\m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net965),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][10] ),
    .A2(net289),
    .B1(net277),
    .B2(\m_blake2.m_hash256.v_q[2][10] ),
    .C1(\m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__and3_2_C_X ),
    .X(\m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_X ));
 sky130_fd_sc_hd__o22a_1 \m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__o22a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_X ),
    .A2(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_X ),
    .B2(net363),
    .X(\m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__o22a_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1099),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][11] ),
    .A2(net294),
    .B1(net405),
    .B2(\m_blake2.m_hash256.v_q[0][11] ),
    .X(\m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net895),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][12] ),
    .A2(net291),
    .B1(net279),
    .B2(\m_blake2.m_hash256.v_q[2][12] ),
    .X(\m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1404),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net301),
    .X(\m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][13] ),
    .A2(net295),
    .B1(\m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__a31o_2_A3_X ),
    .C1(\m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .A2(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_X ),
    .B1(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .Y(\m_blake2.m_hash256.m_g.a0[14]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ),
    .B(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__o32a_4 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X  (.A1(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ),
    .A2(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ),
    .A3(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ),
    .B1(net100),
    .B2(\m_blake2.m_hash256.m_matrix[0][13] ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[6][13] ),
    .A2(net96),
    .B1(net120),
    .B2(\m_blake2.m_hash256.m_matrix[15][13] ),
    .C1(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[13][13] ),
    .A2(net116),
    .B1(net148),
    .B2(\m_blake2.m_hash256.m_matrix[11][13] ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a2111o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[5][13] ),
    .A2(net112),
    .B1(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ),
    .C1(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ),
    .D1(net104),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[4][13] ),
    .A2(net84),
    .B1(net136),
    .B2(\m_blake2.m_hash256.m_matrix[2][13] ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[7][13] ),
    .A2(net108),
    .B1(net132),
    .B2(\m_blake2.m_hash256.m_matrix[3][13] ),
    .C1(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[8][13] ),
    .A2(net128),
    .B1(net144),
    .B2(\m_blake2.m_hash256.m_matrix[10][13] ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[9][13] ),
    .A2(net124),
    .B1(net88),
    .B2(\m_blake2.m_hash256.m_matrix[14][13] ),
    .C1(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X  (.A1(\m_blake2.m_hash256.m_matrix[1][13] ),
    .A2(net140),
    .B1(net92),
    .B2(\m_blake2.m_hash256.m_matrix[12][13] ),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1124),
    .A1(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][14] ),
    .A2(net294),
    .B1(net286),
    .B2(\m_blake2.m_hash256.v_q[3][14] ),
    .X(\m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1136),
    .A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][15] ),
    .A2(net292),
    .B1(net287),
    .B2(\m_blake2.m_hash256.v_q[3][15] ),
    .X(\m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1350),
    .A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][16] ),
    .A2(net289),
    .B1(\m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net362),
    .X(\m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1191),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][17] ),
    .A2(net289),
    .B1(net284),
    .B2(\m_blake2.m_hash256.v_q[3][17] ),
    .X(\m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net922),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][18] ),
    .A2(net289),
    .B1(net285),
    .B2(\m_blake2.m_hash256.v_q[3][18] ),
    .X(\m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1268),
    .A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][19] ),
    .A2(net293),
    .B1(net287),
    .B2(\m_blake2.m_hash256.v_q[3][19] ),
    .X(\m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1192),
    .A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][1] ),
    .A2(net290),
    .B1(net278),
    .B2(\m_blake2.m_hash256.v_q[2][1] ),
    .X(\m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1063),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][20] ),
    .A2(net291),
    .B1(net285),
    .B2(\m_blake2.m_hash256.v_q[3][20] ),
    .X(\m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1108),
    .A1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net301),
    .X(\m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][21] ),
    .A2(net295),
    .B1(net283),
    .B2(\m_blake2.m_hash256.v_q[2][21] ),
    .X(\m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1253),
    .A1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][22] ),
    .A2(net292),
    .B1(net286),
    .B2(\m_blake2.m_hash256.v_q[3][22] ),
    .X(\m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1313),
    .A1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][23] ),
    .A2(net292),
    .B1(net286),
    .B2(\m_blake2.m_hash256.v_q[3][23] ),
    .X(\m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1115),
    .A1(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][24] ),
    .A2(net291),
    .B1(net285),
    .B2(\m_blake2.m_hash256.v_q[3][24] ),
    .X(\m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1226),
    .A1(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net301),
    .X(\m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][25] ),
    .A2(net290),
    .B1(net284),
    .B2(\m_blake2.m_hash256.v_q[3][25] ),
    .X(\m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1002),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][26] ),
    .A2(net289),
    .B1(net285),
    .B2(\m_blake2.m_hash256.v_q[3][26] ),
    .X(\m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1279),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][27] ),
    .A2(net293),
    .B1(net287),
    .B2(\m_blake2.m_hash256.v_q[3][27] ),
    .X(\m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1346),
    .A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][28] ),
    .A2(net295),
    .B1(net283),
    .B2(\m_blake2.m_hash256.v_q[2][28] ),
    .X(\m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1342),
    .A1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][29] ),
    .A2(net294),
    .B1(net286),
    .B2(\m_blake2.m_hash256.v_q[3][29] ),
    .X(\m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1033),
    .A1(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][2] ),
    .A2(net290),
    .B1(net284),
    .B2(\m_blake2.m_hash256.v_q[3][2] ),
    .X(\m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net979),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net301),
    .X(\m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][30] ),
    .A2(net292),
    .B1(net286),
    .B2(\m_blake2.m_hash256.v_q[3][30] ),
    .X(\m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1427),
    .A1(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][31] ),
    .A2(net293),
    .B1(net286),
    .B2(\m_blake2.m_hash256.v_q[3][31] ),
    .X(\m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1234),
    .A1(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][3] ),
    .A2(net293),
    .B1(net281),
    .B2(\m_blake2.m_hash256.v_q[2][3] ),
    .X(\m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1012),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][4] ),
    .A2(net291),
    .B1(net406),
    .B2(\m_blake2.m_hash256.v_q[0][4] ),
    .X(\m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1100),
    .A1(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][5] ),
    .A2(net295),
    .B1(net283),
    .B2(\m_blake2.m_hash256.v_q[2][5] ),
    .X(\m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1196),
    .A1(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net303),
    .X(\m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][6] ),
    .A2(net292),
    .B1(net286),
    .B2(\m_blake2.m_hash256.v_q[3][6] ),
    .X(\m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1312),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][7] ),
    .A2(net293),
    .B1(\m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net390),
    .X(\m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_X ),
    .A2(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .X(\m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1424),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net302),
    .X(\m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][8] ),
    .A2(net290),
    .B1(net278),
    .B2(\m_blake2.m_hash256.v_q[2][8] ),
    .X(\m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1027),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[1][9] ),
    .A2(net289),
    .B1(net277),
    .B2(\m_blake2.m_hash256.v_q[2][9] ),
    .X(\m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[1][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1073),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net300),
    .X(\m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1134),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][0] ),
    .B(\m_blake2.m_hash256.v_q[2][0] ),
    .Y(\m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1369),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][10] ),
    .B(\m_blake2.m_hash256.v_q[2][10] ),
    .Y(\m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][11] ),
    .A2(net282),
    .B1(\m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .Y(\m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net917),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][11] ),
    .B(\m_blake2.m_hash256.v_q[2][11] ),
    .X(\m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1298),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net414),
    .X(\m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][12] ),
    .B(\m_blake2.m_hash256.v_q[2][12] ),
    .Y(\m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][13] ),
    .A2(net283),
    .B1(net406),
    .B2(\m_blake2.m_hash256.v_q[0][13] ),
    .X(\m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1076),
    .A1(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][13] ),
    .B(\m_blake2.m_hash256.v_q[2][13] ),
    .Y(\m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][14] ),
    .A2(net282),
    .B1(\m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net386),
    .X(\m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[2][14] ),
    .A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_2 \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][14] ),
    .B(\m_blake2.m_hash256.v_q[2][14] ),
    .X(\m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][15] ),
    .A2(net280),
    .B1(\m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net389),
    .X(\m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1131),
    .A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][15] ),
    .B(\m_blake2.m_hash256.v_q[2][15] ),
    .X(\m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][16] ),
    .A2(net277),
    .B1(net284),
    .B2(\m_blake2.m_hash256.v_q[3][16] ),
    .X(\m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1774),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][16] ),
    .B(\m_blake2.m_hash256.v_q[2][16] ),
    .X(\m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][17] ),
    .A2(net277),
    .B1(\m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net362),
    .X(\m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1087),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][17] ),
    .B(\m_blake2.m_hash256.v_q[2][17] ),
    .Y(\m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][18] ),
    .A2(net278),
    .B1(\m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net363),
    .X(\m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1649),
    .A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][18] ),
    .B(\m_blake2.m_hash256.v_q[2][18] ),
    .Y(\m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][19] ),
    .A2(net281),
    .B1(\m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net389),
    .X(\m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1168),
    .A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][19] ),
    .B(\m_blake2.m_hash256.v_q[2][19] ),
    .Y(\m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1159),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net414),
    .X(\m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][1] ),
    .B(\m_blake2.m_hash256.v_q[2][1] ),
    .Y(\m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][20] ),
    .A2(net279),
    .B1(\m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net399),
    .X(\m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1008),
    .A1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net414),
    .X(\m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][20] ),
    .B(\m_blake2.m_hash256.v_q[2][20] ),
    .X(\m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1301),
    .A1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][21] ),
    .B(\m_blake2.m_hash256.v_q[2][21] ),
    .Y(\m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][22] ),
    .A2(net282),
    .B1(\m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net386),
    .X(\m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1402),
    .A1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][22] ),
    .B(\m_blake2.m_hash256.v_q[2][22] ),
    .X(\m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][23] ),
    .A2(net280),
    .B1(\m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net389),
    .X(\m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1101),
    .A1(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][23] ),
    .B(\m_blake2.m_hash256.v_q[2][23] ),
    .Y(\m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][24] ),
    .A2(net279),
    .B1(\m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net372),
    .X(\m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1141),
    .A1(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net414),
    .X(\m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][24] ),
    .B(\m_blake2.m_hash256.v_q[2][24] ),
    .Y(\m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][25] ),
    .A2(net278),
    .B1(\m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net366),
    .X(\m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1223),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][25] ),
    .B(\m_blake2.m_hash256.v_q[2][25] ),
    .Y(\m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][26] ),
    .A2(net278),
    .B1(\m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net367),
    .X(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1  (.A1(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .A2(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_X ),
    .B1(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X ),
    .X(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1145),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net414),
    .X(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][26] ),
    .B(\m_blake2.m_hash256.v_q[2][26] ),
    .Y(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__a211oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][27] ),
    .A2(net280),
    .B1(\m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net390),
    .Y(\m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__a211oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1095),
    .A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][27] ),
    .B(\m_blake2.m_hash256.v_q[2][27] ),
    .Y(\m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1396),
    .A1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][28] ),
    .B(\m_blake2.m_hash256.v_q[2][28] ),
    .X(\m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__a211oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][29] ),
    .A2(net283),
    .B1(\m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net379),
    .Y(\m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__a211oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1019),
    .A1(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][29] ),
    .B(\m_blake2.m_hash256.v_q[2][29] ),
    .X(\m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][2] ),
    .A2(net278),
    .B1(net403),
    .B2(\m_blake2.m_hash256.v_q[0][2] ),
    .C1(\m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .X(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_X ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__nor2_2_B  (.A(net367),
    .B(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_X ),
    .Y(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1038),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net414),
    .X(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][2] ),
    .B(\m_blake2.m_hash256.v_q[2][2] ),
    .X(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[74]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][30] ),
    .A2(net280),
    .B1(\m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net389),
    .X(\m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1114),
    .A1(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][30] ),
    .B(\m_blake2.m_hash256.v_q[2][30] ),
    .Y(\m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__a211oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][31] ),
    .A2(net281),
    .B1(\m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net390),
    .Y(\m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__a211oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1197),
    .A1(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][31] ),
    .B(\m_blake2.m_hash256.v_q[2][31] ),
    .Y(\m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1311),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][3] ),
    .B(\m_blake2.m_hash256.v_q[2][3] ),
    .Y(\m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a21oi_1 \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__a21oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][4] ),
    .A2(net279),
    .B1(\m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .Y(\m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1071),
    .A1(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][4] ),
    .B(\m_blake2.m_hash256.v_q[2][4] ),
    .X(\m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1097),
    .A1(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net416),
    .X(\m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][5] ),
    .B(\m_blake2.m_hash256.v_q[2][5] ),
    .Y(\m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][6] ),
    .A2(net282),
    .B1(\m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net387),
    .X(\m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1205),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][6] ),
    .B(\m_blake2.m_hash256.v_q[2][6] ),
    .X(\m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[2][7] ),
    .A2(net280),
    .B1(net287),
    .B2(\m_blake2.m_hash256.v_q[3][7] ),
    .X(\m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1478),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net415),
    .X(\m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][7] ),
    .B(\m_blake2.m_hash256.v_q[2][7] ),
    .Y(\m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1370),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][8] ),
    .B(\m_blake2.m_hash256.v_q[2][8] ),
    .X(\m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[2][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1116),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net413),
    .X(\m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[10][9] ),
    .B(\m_blake2.m_hash256.v_q[2][9] ),
    .Y(\m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[73]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net472),
    .A2(net476),
    .A3(\m_blake2.m_hash256.v_q[3][0] ),
    .B1(net366),
    .X(\m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1153),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][0] ),
    .B(\m_blake2.m_hash256.v_q[3][0] ),
    .Y(\m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__and3_2_C  (.A(net470),
    .B(net475),
    .C(\m_blake2.m_hash256.v_q[3][10] ),
    .X(\m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net968),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][10] ),
    .B(\m_blake2.m_hash256.v_q[3][10] ),
    .Y(\m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net953),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[3][11] ),
    .B(net288),
    .Y(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2  (.A1(net355),
    .A2(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A3(\m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B1(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_B1 ),
    .X(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X ),
    .Y(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][11] ),
    .B(\m_blake2.m_hash256.v_q[3][11] ),
    .Y(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[3][12] ),
    .A2(net285),
    .B1(\m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net372),
    .X(\m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1473),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net418),
    .X(\m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][12] ),
    .B(\m_blake2.m_hash256.v_q[3][12] ),
    .Y(\m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net473),
    .A2(net477),
    .A3(\m_blake2.m_hash256.v_q[3][13] ),
    .B1(net378),
    .X(\m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1323),
    .A1(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][13] ),
    .B(\m_blake2.m_hash256.v_q[3][13] ),
    .Y(\m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1316),
    .A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][14] ),
    .B(\m_blake2.m_hash256.v_q[3][14] ),
    .X(\m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1251),
    .A1(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][15] ),
    .B(\m_blake2.m_hash256.v_q[3][15] ),
    .X(\m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1375),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][16] ),
    .B(\m_blake2.m_hash256.v_q[3][16] ),
    .Y(\m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_70_clk),
    .D(\m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net962),
    .A1(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][17] ),
    .B(\m_blake2.m_hash256.v_q[3][17] ),
    .X(\m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_8_clk),
    .D(\m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net956),
    .A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][18] ),
    .B(\m_blake2.m_hash256.v_q[3][18] ),
    .X(\m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[114]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1327),
    .A1(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][19] ),
    .B(\m_blake2.m_hash256.v_q[3][19] ),
    .Y(\m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[3][1] ),
    .A2(net284),
    .B1(\m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net363),
    .X(\m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1339),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][1] ),
    .B(\m_blake2.m_hash256.v_q[3][1] ),
    .Y(\m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1084),
    .A1(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net418),
    .X(\m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][20] ),
    .B(\m_blake2.m_hash256.v_q[3][20] ),
    .Y(\m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__a211oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[3][21] ),
    .A2(net288),
    .B1(\m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net378),
    .Y(\m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__a211oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1046),
    .A1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][21] ),
    .B(\m_blake2.m_hash256.v_q[3][21] ),
    .Y(\m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1231),
    .A1(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][22] ),
    .B(\m_blake2.m_hash256.v_q[3][22] ),
    .X(\m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[118]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1077),
    .A1(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][23] ),
    .B(\m_blake2.m_hash256.v_q[3][23] ),
    .Y(\m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net976),
    .A1(\m_blake2.m_hash256.m_g.a_q[24]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net418),
    .X(\m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][24] ),
    .B(\m_blake2.m_hash256.v_q[3][24] ),
    .X(\m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1066),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][25] ),
    .B(\m_blake2.m_hash256.v_q[3][25] ),
    .X(\m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1246),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][26] ),
    .B(\m_blake2.m_hash256.v_q[3][26] ),
    .Y(\m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1103),
    .A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][27] ),
    .B(\m_blake2.m_hash256.v_q[3][27] ),
    .Y(\m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[123]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[3][28] ),
    .A2(net288),
    .B1(\m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net378),
    .X(\m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1139),
    .A1(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_A0 ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][28] ),
    .B(\m_blake2.m_hash256.v_q[3][28] ),
    .Y(\m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1162),
    .A1(\m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_X ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][29] ),
    .B(\m_blake2.m_hash256.v_q[3][29] ),
    .X(\m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1389),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net418),
    .X(\m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][2] ),
    .B(\m_blake2.m_hash256.v_q[3][2] ),
    .Y(\m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[98]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1386),
    .A1(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][30] ),
    .B(\m_blake2.m_hash256.v_q[3][30] ),
    .Y(\m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1344),
    .A1(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][31] ),
    .B(\m_blake2.m_hash256.v_q[3][31] ),
    .Y(\m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[135]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[3][3] ),
    .A2(net287),
    .B1(\m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net396),
    .X(\m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1243),
    .A1(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][3] ),
    .B(\m_blake2.m_hash256.v_q[3][3] ),
    .Y(\m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net992),
    .A1(\m_blake2.m_hash256.m_g.a_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_blake2.m_hash256.v_q[3][4] ),
    .B(net288),
    .Y(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2  (.A1(net354),
    .A2(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .A3(\m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .B1(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_B1 ),
    .X(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][4] ),
    .B(\m_blake2.m_hash256.v_q[3][4] ),
    .X(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[100]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_blake2.m_hash256.v_q[3][5] ),
    .A2(net288),
    .B1(\m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net379),
    .X(\m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__a211o_2_A1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1426),
    .A1(\m_blake2.m_hash256.m_g.a_q[5]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net420),
    .X(\m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][5] ),
    .B(\m_blake2.m_hash256.v_q[3][5] ),
    .Y(\m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[109]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1133),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][6] ),
    .B(\m_blake2.m_hash256.v_q[3][6] ),
    .X(\m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1288),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net419),
    .X(\m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][7] ),
    .B(\m_blake2.m_hash256.v_q[3][7] ),
    .Y(\m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[103]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .Y(\m_blake2.m_hash256.h_flat[111]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a211oi_1 \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__a211oi_2_A1  (.A1(\m_blake2.m_hash256.v_q[3][8] ),
    .A2(net284),
    .B1(\m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .C1(net371),
    .Y(\m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__a211oi_2_A1_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1015),
    .A1(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][8] ),
    .B(\m_blake2.m_hash256.v_q[3][8] ),
    .X(\m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a31o_1 \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__a31o_2_A3  (.A1(net472),
    .A2(net476),
    .A3(\m_blake2.m_hash256.v_q[3][9] ),
    .B1(net363),
    .X(\m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__a31o_2_A3_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[3][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net975),
    .A1(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net417),
    .X(\m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__xor2_2_B  (.A(\m_blake2.m_hash256.v_q[11][9] ),
    .B(\m_blake2.m_hash256.v_q[3][9] ),
    .X(\m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[105]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__xor2_2_B_X ),
    .Y(\m_blake2.m_hash256.h_flat[113]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1028),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][0] ),
    .B(\m_blake2.m_hash256.v_q[12][0] ),
    .Y(\m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .B(\m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net928),
    .A1(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][10] ),
    .A1(\m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net370),
    .X(\m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][10] ),
    .B(\m_blake2.m_hash256.v_q[12][10] ),
    .Y(\m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net906),
    .A1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net230),
    .X(\m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][11] ),
    .A1(\m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net375),
    .X(\m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][11] ),
    .B(\m_blake2.m_hash256.v_q[12][11] ),
    .Y(\m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[147]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1652),
    .A1(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][12] ),
    .B(\m_blake2.m_hash256.v_q[12][12] ),
    .Y(\m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net856),
    .A1(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][13] ),
    .A1(\m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net397),
    .X(\m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][13] ),
    .B(\m_blake2.m_hash256.v_q[12][13] ),
    .Y(\m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net930),
    .A1(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][14] ),
    .B(\m_blake2.m_hash256.v_q[12][14] ),
    .Y(\m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net907),
    .A1(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net232),
    .X(\m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][15] ),
    .A1(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net396),
    .X(\m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][15] ),
    .B(\m_blake2.m_hash256.v_q[12][15] ),
    .Y(\m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net934),
    .A1(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net230),
    .X(\m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][16] ),
    .B(\m_blake2.m_hash256.v_q[12][16] ),
    .Y(\m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net901),
    .A1(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][17] ),
    .B(\m_blake2.m_hash256.v_q[12][17] ),
    .Y(\m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net883),
    .A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][18] ),
    .B(\m_blake2.m_hash256.v_q[12][18] ),
    .Y(\m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net886),
    .A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net230),
    .X(\m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][19] ),
    .B(\m_blake2.m_hash256.v_q[12][19] ),
    .Y(\m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1079),
    .A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][1] ),
    .B(\m_blake2.m_hash256.v_q[12][1] ),
    .Y(\m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .B(\m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net936),
    .A1(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][20] ),
    .B(\m_blake2.m_hash256.v_q[12][20] ),
    .Y(\m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[156]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net891),
    .A1(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net232),
    .X(\m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][21] ),
    .A1(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net397),
    .X(\m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][21] ),
    .B(\m_blake2.m_hash256.v_q[12][21] ),
    .Y(\m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[149]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[157]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net959),
    .A1(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][22] ),
    .B(\m_blake2.m_hash256.v_q[12][22] ),
    .Y(\m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net902),
    .A1(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net232),
    .X(\m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][23] ),
    .A1(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net396),
    .X(\m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][23] ),
    .B(\m_blake2.m_hash256.v_q[12][23] ),
    .Y(\m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[151]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[159]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1338),
    .A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][24] ),
    .B(\m_blake2.m_hash256.v_q[12][24] ),
    .Y(\m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net918),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][25] ),
    .A1(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net368),
    .X(\m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][25] ),
    .B(\m_blake2.m_hash256.v_q[12][25] ),
    .Y(\m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net889),
    .A1(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][26] ),
    .A1(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net374),
    .X(\m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][26] ),
    .B(\m_blake2.m_hash256.v_q[12][26] ),
    .Y(\m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net880),
    .A1(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net230),
    .X(\m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[4][27] ),
    .A1(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net375),
    .X(\m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][27] ),
    .B(\m_blake2.m_hash256.v_q[12][27] ),
    .Y(\m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[155]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[4][27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1005),
    .A1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][28] ),
    .B(\m_blake2.m_hash256.v_q[12][28] ),
    .Y(\m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net929),
    .A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net232),
    .X(\m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][29] ),
    .B(\m_blake2.m_hash256.v_q[12][29] ),
    .Y(\m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1872),
    .A1(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.v_q[4][2] ),
    .Y(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][2] ),
    .B(\m_blake2.m_hash256.v_q[12][2] ),
    .Y(\m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net867),
    .A1(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net232),
    .X(\m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][30] ),
    .B(\m_blake2.m_hash256.v_q[12][30] ),
    .Y(\m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net919),
    .A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net232),
    .X(\m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][31] ),
    .B(\m_blake2.m_hash256.v_q[12][31] ),
    .Y(\m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1847),
    .A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__clkinv_2 \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__inv_2_A  (.A(\m_blake2.m_hash256.v_q[4][3] ),
    .Y(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][3] ),
    .B(\m_blake2.m_hash256.v_q[12][3] ),
    .Y(\m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1051),
    .A1(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][4] ),
    .B(\m_blake2.m_hash256.v_q[12][4] ),
    .Y(\m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .B(\m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1181),
    .A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][5] ),
    .B(\m_blake2.m_hash256.v_q[12][5] ),
    .Y(\m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .B(\m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net985),
    .A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net231),
    .X(\m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][6] ),
    .B(\m_blake2.m_hash256.v_q[12][6] ),
    .Y(\m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .B(\m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net869),
    .A1(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net232),
    .X(\m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][7] ),
    .B(\m_blake2.m_hash256.v_q[12][7] ),
    .Y(\m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[143]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net961),
    .A1(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net230),
    .X(\m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][8] ),
    .B(\m_blake2.m_hash256.v_q[12][8] ),
    .Y(\m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[4][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net844),
    .A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net229),
    .X(\m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[4][9] ),
    .B(\m_blake2.m_hash256.v_q[12][9] ),
    .Y(\m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_A1 ),
    .B(\m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][0] ),
    .A2(net188),
    .B1(net195),
    .B2(\m_blake2.m_hash256.v_q[7][0] ),
    .X(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1227),
    .A1(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][0] ),
    .B(\m_blake2.m_hash256.v_q[13][0] ),
    .Y(\m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][10] ),
    .A2(net189),
    .B1(net195),
    .B2(\m_blake2.m_hash256.v_q[7][10] ),
    .X(\m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net343),
    .A2(\m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .C1(net177),
    .X(\m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1215),
    .A1(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][10] ),
    .B(\m_blake2.m_hash256.v_q[13][10] ),
    .X(\m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net877),
    .A1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[5][11] ),
    .A1(\m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net377),
    .X(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1  (.A1(net375),
    .A2(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X ),
    .B2(net188),
    .C1(net178),
    .X(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][11] ),
    .B(\m_blake2.m_hash256.v_q[13][11] ),
    .Y(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][12] ),
    .A2(net192),
    .B1(net200),
    .B2(\m_blake2.m_hash256.v_q[7][12] ),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1142),
    .A1(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][12] ),
    .B(\m_blake2.m_hash256.v_q[13][12] ),
    .Y(\m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][13] ),
    .A2(net191),
    .B1(net200),
    .B2(\m_blake2.m_hash256.v_q[7][13] ),
    .X(\m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net360),
    .A2(\m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ),
    .X(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1102),
    .A1(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][13] ),
    .B(\m_blake2.m_hash256.v_q[13][13] ),
    .Y(\m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][14] ),
    .A2(net190),
    .B1(net198),
    .B2(\m_blake2.m_hash256.v_q[7][14] ),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1239),
    .A1(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net160),
    .X(\m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][14] ),
    .B(\m_blake2.m_hash256.v_q[13][14] ),
    .Y(\m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][15] ),
    .A2(net191),
    .B1(net199),
    .B2(\m_blake2.m_hash256.v_q[7][15] ),
    .X(\m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net359),
    .A2(\m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .C1(net179),
    .X(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1113),
    .A1(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][15] ),
    .B(\m_blake2.m_hash256.v_q[13][15] ),
    .X(\m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][16] ),
    .A2(net188),
    .B1(net196),
    .B2(\m_blake2.m_hash256.v_q[7][16] ),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1391),
    .A1(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net158),
    .X(\m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][16] ),
    .B(\m_blake2.m_hash256.v_q[13][16] ),
    .Y(\m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][17] ),
    .A2(net187),
    .B1(net195),
    .B2(\m_blake2.m_hash256.v_q[7][17] ),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1067),
    .A1(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][17] ),
    .B(\m_blake2.m_hash256.v_q[13][17] ),
    .Y(\m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][18] ),
    .A2(net188),
    .B1(net196),
    .B2(\m_blake2.m_hash256.v_q[7][18] ),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1081),
    .A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][18] ),
    .B(\m_blake2.m_hash256.v_q[13][18] ),
    .Y(\m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][19] ),
    .A2(net188),
    .B1(net196),
    .B2(\m_blake2.m_hash256.v_q[7][19] ),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1152),
    .A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net158),
    .X(\m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][19] ),
    .B(\m_blake2.m_hash256.v_q[13][19] ),
    .Y(\m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[179]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][1] ),
    .A2(net187),
    .B1(net195),
    .B2(\m_blake2.m_hash256.v_q[7][1] ),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1001),
    .A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][1] ),
    .B(\m_blake2.m_hash256.v_q[13][1] ),
    .Y(\m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][20] ),
    .A2(net192),
    .B1(net200),
    .B2(\m_blake2.m_hash256.v_q[7][20] ),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1106),
    .A1(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][20] ),
    .B(\m_blake2.m_hash256.v_q[13][20] ),
    .Y(\m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][21] ),
    .A2(net191),
    .B1(net199),
    .B2(\m_blake2.m_hash256.v_q[7][21] ),
    .X(\m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net360),
    .A2(\m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .C1(net179),
    .X(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1061),
    .A1(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net160),
    .X(\m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][21] ),
    .B(\m_blake2.m_hash256.v_q[13][21] ),
    .X(\m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[181]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][22] ),
    .A2(net192),
    .B1(net198),
    .B2(\m_blake2.m_hash256.v_q[7][22] ),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1183),
    .A1(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net160),
    .X(\m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][22] ),
    .B(\m_blake2.m_hash256.v_q[13][22] ),
    .X(\m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][23] ),
    .A2(net191),
    .B1(net199),
    .B2(\m_blake2.m_hash256.v_q[7][23] ),
    .X(\m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net359),
    .A2(\m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .C1(net180),
    .X(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1009),
    .A1(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][23] ),
    .B(\m_blake2.m_hash256.v_q[13][23] ),
    .X(\m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[183]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][24] ),
    .A2(net190),
    .B1(net198),
    .B2(\m_blake2.m_hash256.v_q[7][24] ),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_31_clk),
    .D(\m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1180),
    .A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net160),
    .X(\m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][24] ),
    .B(\m_blake2.m_hash256.v_q[13][24] ),
    .Y(\m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[184]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][25] ),
    .A2(net187),
    .B1(net195),
    .B2(\m_blake2.m_hash256.v_q[7][25] ),
    .X(\m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net343),
    .A2(\m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ),
    .X(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net932),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][25] ),
    .B(\m_blake2.m_hash256.v_q[13][25] ),
    .Y(\m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][26] ),
    .A2(net189),
    .B1(net197),
    .B2(\m_blake2.m_hash256.v_q[7][26] ),
    .X(\m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a211o_1 \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2  (.A1(net348),
    .A2(\m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ),
    .C1(net177),
    .X(\m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1434),
    .A1(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][26] ),
    .B(\m_blake2.m_hash256.v_q[13][26] ),
    .X(\m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][27] ),
    .A2(net189),
    .B1(net197),
    .B2(\m_blake2.m_hash256.v_q[7][27] ),
    .X(\m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net350),
    .A2(\m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ),
    .X(\m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1075),
    .A1(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net158),
    .X(\m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][27] ),
    .B(\m_blake2.m_hash256.v_q[13][27] ),
    .Y(\m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[187]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][28] ),
    .A2(net190),
    .B1(net198),
    .B2(\m_blake2.m_hash256.v_q[7][28] ),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net977),
    .A1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net160),
    .X(\m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][28] ),
    .B(\m_blake2.m_hash256.v_q[13][28] ),
    .Y(\m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][29] ),
    .A2(net191),
    .B1(net199),
    .B2(\m_blake2.m_hash256.v_q[7][29] ),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1041),
    .A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][29] ),
    .B(\m_blake2.m_hash256.v_q[13][29] ),
    .X(\m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[189]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][2] ),
    .A2(net187),
    .B1(net195),
    .B2(\m_blake2.m_hash256.v_q[7][2] ),
    .X(\m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net978),
    .A1(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][2] ),
    .B(\m_blake2.m_hash256.v_q[13][2] ),
    .Y(\m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][30] ),
    .A2(net192),
    .B1(net200),
    .B2(\m_blake2.m_hash256.v_q[7][30] ),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1185),
    .A1(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][30] ),
    .B(\m_blake2.m_hash256.v_q[13][30] ),
    .Y(\m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net937),
    .A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__mux2_1_A0_1  (.A0(\m_blake2.m_hash256.v_q[5][31] ),
    .A1(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net396),
    .X(\m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__mux2_1_A0_1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][31] ),
    .B(\m_blake2.m_hash256.v_q[13][31] ),
    .Y(\m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[191]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][3] ),
    .A2(net190),
    .B1(net198),
    .B2(\m_blake2.m_hash256.v_q[7][3] ),
    .X(\m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1020),
    .A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net158),
    .X(\m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][3] ),
    .B(\m_blake2.m_hash256.v_q[13][3] ),
    .Y(\m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][4] ),
    .A2(net190),
    .B1(net198),
    .B2(\m_blake2.m_hash256.v_q[7][4] ),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net971),
    .A1(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net160),
    .X(\m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][4] ),
    .B(\m_blake2.m_hash256.v_q[13][4] ),
    .Y(\m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][5] ),
    .A2(net192),
    .B1(net200),
    .B2(\m_blake2.m_hash256.v_q[7][5] ),
    .X(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net972),
    .A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][5] ),
    .B(\m_blake2.m_hash256.v_q[13][5] ),
    .Y(\m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[165]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][6] ),
    .A2(net190),
    .B1(net198),
    .B2(\m_blake2.m_hash256.v_q[7][6] ),
    .X(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1258),
    .A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net160),
    .X(\m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][6] ),
    .B(\m_blake2.m_hash256.v_q[13][6] ),
    .Y(\m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][7] ),
    .A2(net191),
    .B1(net199),
    .B2(\m_blake2.m_hash256.v_q[7][7] ),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1308),
    .A1(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net159),
    .X(\m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][7] ),
    .B(\m_blake2.m_hash256.v_q[13][7] ),
    .X(\m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[167]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][8] ),
    .A2(net189),
    .B1(net196),
    .B2(\m_blake2.m_hash256.v_q[7][8] ),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1617),
    .A1(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net158),
    .X(\m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][8] ),
    .B(\m_blake2.m_hash256.v_q[13][8] ),
    .X(\m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[168]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[5][9] ),
    .A2(net187),
    .B1(net195),
    .B2(\m_blake2.m_hash256.v_q[7][9] ),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[5][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1054),
    .A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net157),
    .X(\m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[5][9] ),
    .B(\m_blake2.m_hash256.v_q[13][9] ),
    .Y(\m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_29_clk),
    .D(\m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net948),
    .S(net216),
    .X(\m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][0] ),
    .A1(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net374),
    .X(\m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][0] ),
    .B(\m_blake2.m_hash256.v_q[14][0] ),
    .Y(\m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[192]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][10] ),
    .A1(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net370),
    .X(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(net344),
    .A2_N(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net255),
    .X(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net957),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][10] ),
    .B(\m_blake2.m_hash256.v_q[14][10] ),
    .Y(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[6][11] ),
    .A2(net256),
    .B1(net196),
    .B2(\m_blake2.m_hash256.v_q[7][11] ),
    .X(\m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1_X ));
 sky130_fd_sc_hd__a21o_1 \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2  (.A1(net349),
    .A2(\m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1_X ),
    .B1(\m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1_X ),
    .X(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1160),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][11] ),
    .B(\m_blake2.m_hash256.v_q[14][11] ),
    .Y(\m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][12] ),
    .A1(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net395),
    .X(\m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1039),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][12] ),
    .B(\m_blake2.m_hash256.v_q[14][12] ),
    .Y(\m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][13] ),
    .A1(\m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net397),
    .X(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2  (.A1(net257),
    .A2(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X ),
    .B2(net397),
    .C1(net179),
    .X(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1037),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][13] ),
    .B(\m_blake2.m_hash256.v_q[14][13] ),
    .Y(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][14] ),
    .A1(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net380),
    .X(\m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1107),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][14] ),
    .B(\m_blake2.m_hash256.v_q[14][14] ),
    .Y(\m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][15] ),
    .A1(\m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net396),
    .X(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(net359),
    .A2_N(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net257),
    .X(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1203),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][15] ),
    .B(\m_blake2.m_hash256.v_q[14][15] ),
    .Y(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][16] ),
    .A1(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net380),
    .X(\m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1055),
    .S(net216),
    .X(\m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][16] ),
    .B(\m_blake2.m_hash256.v_q[14][16] ),
    .Y(\m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][17] ),
    .A1(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net367),
    .X(\m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1034),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][17] ),
    .B(\m_blake2.m_hash256.v_q[14][17] ),
    .Y(\m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][18] ),
    .A1(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net373),
    .X(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net939),
    .S(net216),
    .X(\m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][18] ),
    .B(\m_blake2.m_hash256.v_q[14][18] ),
    .Y(\m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][19] ),
    .A1(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net375),
    .X(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1409),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][19] ),
    .B(\m_blake2.m_hash256.v_q[14][19] ),
    .Y(\m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net905),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][1] ),
    .A1(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net371),
    .X(\m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][1] ),
    .B(\m_blake2.m_hash256.v_q[14][1] ),
    .Y(\m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][20] ),
    .A1(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net395),
    .X(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1219),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][20] ),
    .B(\m_blake2.m_hash256.v_q[14][20] ),
    .Y(\m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][21] ),
    .A1(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net397),
    .X(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(net360),
    .A2_N(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net257),
    .X(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net931),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][21] ),
    .B(\m_blake2.m_hash256.v_q[14][21] ),
    .Y(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[213]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][22] ),
    .A1(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net383),
    .X(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net933),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][22] ),
    .B(\m_blake2.m_hash256.v_q[14][22] ),
    .Y(\m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][23] ),
    .A1(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net397),
    .X(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(net360),
    .A2_N(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_X ),
    .B1(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net257),
    .X(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1089),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][23] ),
    .B(\m_blake2.m_hash256.v_q[14][23] ),
    .Y(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[215]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][24] ),
    .A1(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net380),
    .X(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1110),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][24] ),
    .B(\m_blake2.m_hash256.v_q[14][24] ),
    .Y(\m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][25] ),
    .A1(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net368),
    .X(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2  (.A1(net255),
    .A2(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .B2(net368),
    .C1(net177),
    .X(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1031),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][25] ),
    .B(\m_blake2.m_hash256.v_q[14][25] ),
    .Y(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][26] ),
    .A1(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net369),
    .X(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a2bb2o_1 \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1  (.A1_N(net348),
    .A2_N(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_X ),
    .B1(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B2(net255),
    .X(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net982),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][26] ),
    .B(\m_blake2.m_hash256.v_q[14][26] ),
    .Y(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][27] ),
    .A1(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net375),
    .X(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2  (.A1(net256),
    .A2(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X ),
    .B1(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_X ),
    .B2(net375),
    .C1(net178),
    .X(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_X ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net955),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][27] ),
    .B(\m_blake2.m_hash256.v_q[14][27] ),
    .Y(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[219]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][28] ),
    .A1(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net384),
    .X(\m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1463),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][28] ),
    .B(\m_blake2.m_hash256.v_q[14][28] ),
    .Y(\m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][29] ),
    .A1(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net397),
    .X(\m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1204),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][29] ),
    .B(\m_blake2.m_hash256.v_q[14][29] ),
    .Y(\m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1036),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][2] ),
    .A1(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net369),
    .X(\m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][2] ),
    .B(\m_blake2.m_hash256.v_q[14][2] ),
    .Y(\m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][30] ),
    .A1(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net392),
    .X(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net944),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][30] ),
    .B(\m_blake2.m_hash256.v_q[14][30] ),
    .Y(\m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[6][31] ),
    .A2(net258),
    .B1(net199),
    .B2(\m_blake2.m_hash256.v_q[7][31] ),
    .X(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1591),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][31] ),
    .B(\m_blake2.m_hash256.v_q[14][31] ),
    .Y(\m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net921),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][3] ),
    .A1(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net381),
    .X(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][3] ),
    .B(\m_blake2.m_hash256.v_q[14][3] ),
    .Y(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net951),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][4] ),
    .A1(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net384),
    .X(\m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][4] ),
    .B(\m_blake2.m_hash256.v_q[14][4] ),
    .Y(\m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[196]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net945),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][5] ),
    .A1(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net397),
    .X(\m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][5] ),
    .B(\m_blake2.m_hash256.v_q[14][5] ),
    .Y(\m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[197]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net987),
    .S(net214),
    .X(\m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][6] ),
    .A1(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net383),
    .X(\m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][6] ),
    .B(\m_blake2.m_hash256.v_q[14][6] ),
    .Y(\m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1030),
    .S(net215),
    .X(\m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][7] ),
    .A1(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net396),
    .X(\m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][7] ),
    .B(\m_blake2.m_hash256.v_q[14][7] ),
    .Y(\m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[199]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1062),
    .S(net216),
    .X(\m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][8] ),
    .A1(\m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__or2_2_B_X ),
    .S(net376),
    .X(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][8] ),
    .B(\m_blake2.m_hash256.v_q[14][8] ),
    .Y(\m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[6][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1074),
    .S(net213),
    .X(\m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[6][9] ),
    .A1(\m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net367),
    .X(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[6][9] ),
    .B(\m_blake2.m_hash256.v_q[14][9] ),
    .Y(\m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1280),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][0] ),
    .B(\m_blake2.m_hash256.v_q[15][0] ),
    .Y(\m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1505),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][10] ),
    .B(\m_blake2.m_hash256.v_q[15][10] ),
    .X(\m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1228),
    .S(net204),
    .X(\m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][11] ),
    .B(\m_blake2.m_hash256.v_q[15][11] ),
    .X(\m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1459),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][12] ),
    .B(\m_blake2.m_hash256.v_q[15][12] ),
    .Y(\m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1471),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][13] ),
    .B(\m_blake2.m_hash256.v_q[15][13] ),
    .Y(\m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1523),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][14] ),
    .B(\m_blake2.m_hash256.v_q[15][14] ),
    .Y(\m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1792),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][15] ),
    .B(\m_blake2.m_hash256.v_q[15][15] ),
    .X(\m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_48_clk),
    .D(\m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1510),
    .S(net204),
    .X(\m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][16] ),
    .B(\m_blake2.m_hash256.v_q[15][16] ),
    .Y(\m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1495),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][17] ),
    .B(\m_blake2.m_hash256.v_q[15][17] ),
    .Y(\m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1202),
    .S(net204),
    .X(\m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][18] ),
    .B(\m_blake2.m_hash256.v_q[15][18] ),
    .Y(\m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1439),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][19] ),
    .B(\m_blake2.m_hash256.v_q[15][19] ),
    .Y(\m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[243]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1229),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][1] ),
    .B(\m_blake2.m_hash256.v_q[15][1] ),
    .X(\m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1490),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][20] ),
    .B(\m_blake2.m_hash256.v_q[15][20] ),
    .Y(\m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_40_clk),
    .D(\m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1390),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][21] ),
    .B(\m_blake2.m_hash256.v_q[15][21] ),
    .X(\m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1222),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][22] ),
    .B(\m_blake2.m_hash256.v_q[15][22] ),
    .X(\m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1423),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][23] ),
    .B(\m_blake2.m_hash256.v_q[15][23] ),
    .X(\m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1704),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][24] ),
    .B(\m_blake2.m_hash256.v_q[15][24] ),
    .Y(\m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__a22o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1607),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][25] ),
    .B(\m_blake2.m_hash256.v_q[15][25] ),
    .Y(\m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__a22o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1436),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][26] ),
    .B(\m_blake2.m_hash256.v_q[15][26] ),
    .Y(\m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__a22o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1245),
    .S(net204),
    .X(\m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][27] ),
    .B(\m_blake2.m_hash256.v_q[15][27] ),
    .Y(\m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__a22o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_35_clk),
    .D(\m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1599),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][28] ),
    .B(\m_blake2.m_hash256.v_q[15][28] ),
    .Y(\m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__a22o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_39_clk),
    .D(\m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1557),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][29] ),
    .B(\m_blake2.m_hash256.v_q[15][29] ),
    .Y(\m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__a22o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1497),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][2] ),
    .B(\m_blake2.m_hash256.v_q[15][2] ),
    .Y(\m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1262),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][30] ),
    .B(\m_blake2.m_hash256.v_q[15][30] ),
    .X(\m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__a22o_2_A1_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1347),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][31] ),
    .B(\m_blake2.m_hash256.v_q[15][31] ),
    .X(\m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B  (.A(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__a32o_2_B1_A3 ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B  (.A(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__xor2_2_A_X ),
    .X(\m_blake2.m_hash256.h_flat[255]_sky130_fd_sc_hd__a32o_2_B1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_36_clk),
    .D(\m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1130),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][3] ),
    .B(\m_blake2.m_hash256.v_q[15][3] ),
    .Y(\m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1305),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][4] ),
    .B(\m_blake2.m_hash256.v_q[15][4] ),
    .Y(\m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1123),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][5] ),
    .B(\m_blake2.m_hash256.v_q[15][5] ),
    .X(\m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[229]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[237]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1190),
    .S(net203),
    .X(\m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][6] ),
    .B(\m_blake2.m_hash256.v_q[15][6] ),
    .Y(\m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1296),
    .S(net202),
    .X(\m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][7] ),
    .B(\m_blake2.m_hash256.v_q[15][7] ),
    .Y(\m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[231]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1440),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][8] ),
    .B(\m_blake2.m_hash256.v_q[15][8] ),
    .X(\m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[240]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[7][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1431),
    .S(net201),
    .X(\m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[7][9] ),
    .B(\m_blake2.m_hash256.v_q[15][9] ),
    .Y(\m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1601),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[8][0] ),
    .A2(net366),
    .B1(net254),
    .X(\m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.v_q[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][10]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .A1(net1345),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[8][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][11]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1361),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[8][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][12]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .A1(net1428),
    .S(net222),
    .X(\m_blake2.m_hash256.v_q[8][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[8][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][13]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1317),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[8][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][14]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1670),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[8][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][15]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1422),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[8][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][16]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .A1(net1838),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[8][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][17]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(\m_blake2.m_hash256.v_q[8][17] ),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_65_clk),
    .D(\m_blake2.m_hash256.v_q[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][18]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .A1(net1472),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[8][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][19]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1536),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1851),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .A1(net1462),
    .S(net222),
    .X(\m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux4_1 \m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__mux4_2_A0  (.A0(\m_blake2.m_hash256.v_q[8][20] ),
    .A1(\m_blake2.m_hash256.v_q[9][20] ),
    .A2(\m_blake2.m_hash256.v_q[10][20] ),
    .A3(\m_blake2.m_hash256.v_q[11][20] ),
    .S0(net477),
    .S1(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ),
    .X(\m_blake2.m_hash256.g_c_buf[20]_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[8][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][21]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1232),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[8][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][22]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1454),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[8][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][23]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1865),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[8][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][24]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .A1(net1470),
    .S(net222),
    .X(\m_blake2.m_hash256.v_q[8][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1394),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[8][25] ),
    .B(net175),
    .X(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__nand2_1 \m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(net355),
    .B(net253),
    .Y(\m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][26]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(net1576),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[8][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][27]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1826),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[8][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][28]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1586),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[8][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][29]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1469),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1855),
    .S(net222),
    .X(\m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[8][2] ),
    .A2(net370),
    .B1(net254),
    .X(\m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[8][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][30]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1210),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[8][30]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[8][30] ),
    .B(net387),
    .X(\m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.v_q[8][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][31]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1726),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[8][3] ),
    .A2(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ),
    .B1(\m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net173),
    .X(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_B1 ));
 sky130_fd_sc_hd__and2_2 \m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2_sky130_fd_sc_hd__and2_2_X  (.A(net355),
    .B(net253),
    .X(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_45_clk),
    .D(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1410),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .A1(net1606),
    .S(net224),
    .X(\m_blake2.m_hash256.v_q[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .A1(net1479),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1398),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[8][6]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[8][6] ),
    .A2(net386),
    .B1(net253),
    .X(\m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[8][7] ),
    .A2(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ),
    .B1(\m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__or2_2_A_X ),
    .B2(net252),
    .X(\m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_54_clk),
    .D(\m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .A1(net1514),
    .S(net223),
    .X(\m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .A1(net1365),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[8][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[8][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .A1(\m_blake2.m_hash256.v_q[8][9] ),
    .S(net221),
    .X(\m_blake2.m_hash256.v_q[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][0] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1378),
    .A1(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][0] ),
    .A2(net366),
    .B1(net250),
    .X(\m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][0] ),
    .B(\m_blake2.m_hash256.v_q[1][0] ),
    .Y(\m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_9_clk),
    .D(\m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][10] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1722),
    .A1(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][10] ),
    .A2(net363),
    .B1(net250),
    .X(\m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][10] ),
    .B(\m_blake2.m_hash256.v_q[1][10] ),
    .Y(\m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_51_clk),
    .D(\m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][11] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1494),
    .A1(\m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and3_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21ai_1 \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][11] ),
    .A2(net388),
    .B1(net249),
    .Y(\m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][11] ),
    .B(\m_blake2.m_hash256.v_q[1][11] ),
    .X(\m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__a32o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][12] ),
    .A2(net350),
    .A3(net252),
    .B1(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B2(\m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][12] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1117),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .S(net154),
    .X(\m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][12] ),
    .B(\m_blake2.m_hash256.v_q[1][12] ),
    .Y(\m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][13] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1522),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][13] ),
    .A2(net379),
    .B1(net251),
    .X(\m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][13] ),
    .B(\m_blake2.m_hash256.v_q[1][13] ),
    .Y(\m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a311o_1 \m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__a311o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][14] ),
    .A2(net354),
    .A3(net249),
    .B1(\m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .C1(\m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.g_c_buf[14]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][14] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1539),
    .A1(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][14] ),
    .B(\m_blake2.m_hash256.v_q[1][14] ),
    .Y(\m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_56_clk),
    .D(\m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][15] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[9][15] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][15] ),
    .A2(net386),
    .B1(net251),
    .X(\m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_A3 ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][15] ),
    .B(\m_blake2.m_hash256.v_q[1][15] ),
    .X(\m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][16] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1356),
    .A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][16] ),
    .A2(net365),
    .B1(net250),
    .X(\m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__o21a_2_A1_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][16] ),
    .B(\m_blake2.m_hash256.v_q[1][16] ),
    .Y(\m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_69_clk),
    .D(\m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][17] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1679),
    .A1(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][17] ),
    .A2(net365),
    .B1(net250),
    .X(\m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_C1 ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][17] ),
    .B(\m_blake2.m_hash256.v_q[1][17] ),
    .X(\m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][18] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[9][18] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][18] ),
    .A2(net364),
    .B1(net250),
    .X(\m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_B1 ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][18] ),
    .B(\m_blake2.m_hash256.v_q[1][18] ),
    .X(\m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a311o_1 \m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__a311o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][19] ),
    .A2(net355),
    .A3(net249),
    .B1(\m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .C1(\m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__o21a_2_A1_X ),
    .X(\m_blake2.m_hash256.g_c_buf[19]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][19] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1764),
    .A1(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][19] ),
    .B(\m_blake2.m_hash256.v_q[1][19] ),
    .Y(\m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[51]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__a32o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][1] ),
    .A2(net346),
    .A3(net249),
    .B1(net169),
    .B2(\m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_66_clk),
    .D(\m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][1] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1753),
    .A1(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][1] ),
    .B(\m_blake2.m_hash256.v_q[1][1] ),
    .Y(\m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_62_clk),
    .D(\m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][20] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net927),
    .A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net154),
    .X(\m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][20] ),
    .B(\m_blake2.m_hash256.v_q[1][20] ),
    .X(\m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][21] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1053),
    .A1(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[9][21] ),
    .B(net379),
    .X(\m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][21] ),
    .B(\m_blake2.m_hash256.v_q[1][21] ),
    .Y(\m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_58_clk),
    .D(\m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][22] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1648),
    .A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][22] ),
    .A2(net387),
    .B1(net251),
    .X(\m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_D1 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][22] ),
    .B(\m_blake2.m_hash256.v_q[1][22] ),
    .Y(\m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[54]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__a22o_2_B1  (.A1(net408),
    .A2(\m_blake2.m_hash256.v_q[10][23] ),
    .B1(\m_blake2.m_hash256.v_q[9][23] ),
    .B2(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ),
    .X(\m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][23] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[9][23] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][23] ),
    .B(\m_blake2.m_hash256.v_q[1][23] ),
    .Y(\m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_61_clk),
    .D(\m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][24] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net897),
    .A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2_2_B_X ),
    .S(net154),
    .X(\m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[9][24] ),
    .B(net372),
    .X(\m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][24] ),
    .B(\m_blake2.m_hash256.v_q[1][24] ),
    .X(\m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][25] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1098),
    .A1(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or3_1 \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B  (.A(net407),
    .B(\m_blake2.m_hash256.v_q[9][25] ),
    .C(net366),
    .X(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_X ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][25] ),
    .B(\m_blake2.m_hash256.v_q[1][25] ),
    .X(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__a32o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][26] ),
    .A2(net345),
    .A3(net250),
    .B1(net171),
    .B2(\m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][26] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[9][26] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][26] ),
    .B(\m_blake2.m_hash256.v_q[1][26] ),
    .Y(\m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[58]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[66]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_52_clk),
    .D(\m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][27] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_blake2.m_hash256.v_q[9][27] ),
    .A1(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o31a_1 \m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__o31a_2_A2  (.A1(net408),
    .A2(\m_blake2.m_hash256.v_q[9][27] ),
    .A3(net388),
    .B1(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ),
    .X(\m_blake2.m_hash256.g_c_buf[27]_sky130_fd_sc_hd__o22a_2_X_B2 ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][27] ),
    .B(\m_blake2.m_hash256.v_q[1][27] ),
    .Y(\m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[59]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_60_clk),
    .D(\m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][28] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net940),
    .A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[9][28] ),
    .B(net378),
    .X(\m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][28] ),
    .B(\m_blake2.m_hash256.v_q[1][28] ),
    .X(\m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][29] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1309),
    .A1(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][29] ),
    .A2(net386),
    .B1(net251),
    .X(\m_blake2.m_hash256.g_c_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2 ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][29] ),
    .B(\m_blake2.m_hash256.v_q[1][29] ),
    .X(\m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][2] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1773),
    .A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net154),
    .X(\m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__o21a_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][2] ),
    .A2(net370),
    .B1(net250),
    .X(\m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][2] ),
    .B(\m_blake2.m_hash256.v_q[1][2] ),
    .X(\m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a221o_1 \m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__a221o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][30] ),
    .A2(net251),
    .B1(net172),
    .B2(\m_blake2.m_hash256.v_q[11][30] ),
    .C1(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(\m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_57_clk),
    .D(\m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][30] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1672),
    .A1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][30] ),
    .B(\m_blake2.m_hash256.v_q[1][30] ),
    .Y(\m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][31] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__mux2_1_A0  (.A0(net1863),
    .A1(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_X_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[9][31] ),
    .B(net388),
    .X(\m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][31] ),
    .B(\m_blake2.m_hash256.v_q[1][31] ),
    .Y(\m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[63]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][3] ),
    .A2(net251),
    .B1(net170),
    .B2(\m_blake2.m_hash256.v_q[10][3] ),
    .X(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_44_clk),
    .D(\m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][3] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1724),
    .A1(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][3] ),
    .B(\m_blake2.m_hash256.v_q[1][3] ),
    .Y(\m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[35]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__a32o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][4] ),
    .A2(net354),
    .A3(net251),
    .B1(net170),
    .B2(\m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][4] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1540),
    .A1(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][4] ),
    .B(\m_blake2.m_hash256.v_q[1][4] ),
    .Y(\m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__and3_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A  (.A(\m_blake2.m_hash256.v_q[9][5] ),
    .B(net354),
    .C(net249),
    .X(\m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_A1 ));
 sky130_fd_sc_hd__nor2_2 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B  (.A(net408),
    .B(net249),
    .Y(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1  (.A(net477),
    .B(net249),
    .Y(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_Y ));
 sky130_fd_sc_hd__or2_4 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_A ),
    .B(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__and2_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_A_sky130_fd_sc_hd__and2_2_X  (.A(net466),
    .B(net469),
    .X(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_A ));
 sky130_fd_sc_hd__nor2_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nor2_2_Y  (.A(net466),
    .B(net469),
    .Y(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_59_clk),
    .D(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][5] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1214),
    .A1(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][5] ),
    .B(\m_blake2.m_hash256.v_q[1][5] ),
    .Y(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a22o_1 \m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__a22o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][6] ),
    .A2(net251),
    .B1(net172),
    .B2(\m_blake2.m_hash256.v_q[11][6] ),
    .X(\m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_55_clk),
    .D(\m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][6] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1634),
    .A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net155),
    .X(\m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][6] ),
    .B(\m_blake2.m_hash256.v_q[1][6] ),
    .Y(\m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_53_clk),
    .D(\m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][7] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1721),
    .A1(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .S(net156),
    .X(\m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[9][7] ),
    .B(net388),
    .X(\m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][7] ),
    .B(\m_blake2.m_hash256.v_q[1][7] ),
    .Y(\m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__a32o_1 \m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__a32o_2_A1  (.A1(\m_blake2.m_hash256.v_q[9][8] ),
    .A2(net346),
    .A3(net250),
    .B1(net171),
    .B2(\m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__or2_2_A_X ),
    .X(\m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_68_clk),
    .D(\m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][8] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1329),
    .A1(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][8] ),
    .B(\m_blake2.m_hash256.v_q[1][8] ),
    .Y(\m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X ),
    .B(\m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_67_clk),
    .D(\m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_blake2.m_hash256.v_q[9][9] ));
 sky130_fd_sc_hd__mux2_1 \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X  (.A0(net1882),
    .A1(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ),
    .S(net153),
    .X(\m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__or2_2_A  (.A(\m_blake2.m_hash256.v_q[9][9] ),
    .B(net362),
    .X(\m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__xor2_1 \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_blake2.m_hash256.v_q[9][9] ),
    .B(\m_blake2.m_hash256.v_q[1][9] ),
    .X(\m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__xnor2_1 \m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B  (.A(\m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .B(\m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.cmd[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.cmd[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.cmd[1] ));
 sky130_fd_sc_hd__and3_1 \m_io.cmd[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net12),
    .X(\m_io.cmd[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.cmd[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.cmd[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.cmd[2] ));
 sky130_fd_sc_hd__and3_1 \m_io.cmd[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net13),
    .X(\m_io.cmd[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nor2_1 \m_io.cmd[2]_sky130_fd_sc_hd__nor2_2_A  (.A(\m_io.cmd[2] ),
    .B(\m_io.cmd[1] ),
    .Y(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__o21ai_2 \m_io.cmd[2]_sky130_fd_sc_hd__o21ai_2_A1  (.A1(\m_io.cmd[2] ),
    .A2(\m_io.cmd[1] ),
    .B1(\m_io.m_config.valid_i ),
    .Y(\m_io.cmd[2]_sky130_fd_sc_hd__o21ai_2_A1_Y ));
 sky130_fd_sc_hd__and2b_2 \m_io.cmd[4]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_io.cmd[5] ),
    .B(\m_io.cmd[4] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2));
 sky130_fd_sc_hd__dfxtp_1 \m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.cmd[4] ));
 sky130_fd_sc_hd__and2_1 \m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X  (.A(net610),
    .B(\m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.cmd[4] ),
    .A1(net14),
    .S(\m_io.en_q ),
    .X(\m_io.cmd[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__and2b_1 \m_io.cmd[5]_sky130_fd_sc_hd__and2b_2_B  (.A_N(\m_io.cmd[4] ),
    .B(\m_io.cmd[5] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2));
 sky130_fd_sc_hd__dfxtp_1 \m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.cmd[5] ));
 sky130_fd_sc_hd__and2_1 \m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X  (.A(net615),
    .B(\m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B ),
    .X(\m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__mux2_1_X  (.A0(\m_io.cmd[5] ),
    .A1(net15),
    .S(\m_io.en_q ),
    .X(\m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_B ));
 sky130_fd_sc_hd__a21oi_1 \m_io.data_v_early_sky130_fd_sc_hd__a21oi_2_A2  (.A1(\m_io.m_block_data.data_cnt_q[0] ),
    .A2(\m_io.data_v_early ),
    .B1(net636),
    .Y(\m_io.data_v_early_sky130_fd_sc_hd__a21oi_2_A2_Y ));
 sky130_fd_sc_hd__and3_1 \m_io.data_v_early_sky130_fd_sc_hd__and3_2_C  (.A(\m_io.m_block_data.data_cnt_q[1] ),
    .B(\m_io.m_block_data.data_cnt_q[0] ),
    .C(\m_io.data_v_early ),
    .X(\m_io.data_v_early_sky130_fd_sc_hd__and3_2_C_X ));
 sky130_fd_sc_hd__inv_2 \m_io.data_v_early_sky130_fd_sc_hd__inv_2_Y  (.A(net308),
    .Y(\m_io.data_v_early ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.en_q_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.en_q_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.en_q ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.hash_v_o_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_19_clk),
    .D(hash_v),
    .Q(\m_io.hash_v_o ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_block_data.data_cnt_q[0] ));
 sky130_fd_sc_hd__nor2_1 \m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(ena_sky130_fd_sc_hd__or2_2_B_A),
    .B(\m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__mux2_1_X  (.A0(net308),
    .A1(\m_io.m_config.valid_i ),
    .S(\m_io.m_block_data.data_cnt_q[0] ),
    .X(\m_io.m_block_data.data_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_block_data.data_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_block_data.data_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_block_data.data_cnt_q[1] ));
 sky130_fd_sc_hd__nor3_1 \m_io.m_block_data.data_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y  (.A(\m_io.data_v_early_sky130_fd_sc_hd__and3_2_C_X ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y ),
    .C(\m_io.data_v_early_sky130_fd_sc_hd__a21oi_2_A2_Y ),
    .Y(\m_io.m_block_data.data_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_block_data.data_cnt_q[2] ));
 sky130_fd_sc_hd__o21a_1 \m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_io.m_block_data.data_cnt_q[2] ),
    .A2(\m_io.data_v_early_sky130_fd_sc_hd__and3_2_C_X ),
    .B1(\m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_block_data.data_cnt_q[2] ),
    .A2(\m_io.data_v_early_sky130_fd_sc_hd__and3_2_C_X ),
    .B1(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y ),
    .Y(\m_io.m_block_data.data_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_block_data.data_cnt_q[3] ));
 sky130_fd_sc_hd__nor3_1 \m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y  (.A(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_B ),
    .C(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_C ),
    .Y(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21oi_1 \m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y  (.A1(\m_io.m_block_data.data_cnt_q[2] ),
    .A2(\m_io.data_v_early_sky130_fd_sc_hd__and3_2_C_X ),
    .B1(net637),
    .Y(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_B ));
 sky130_fd_sc_hd__and3_1 \m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__and3_2_X  (.A(\m_io.m_block_data.data_cnt_q[3] ),
    .B(\m_io.m_block_data.data_cnt_q[2] ),
    .C(\m_io.data_v_early_sky130_fd_sc_hd__and3_2_C_X ),
    .X(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_block_data.data_cnt_q[4] ));
 sky130_fd_sc_hd__and3b_1 \m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B ),
    .C(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_io.m_block_data.data_cnt_q[4] ),
    .B(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_C ),
    .X(\m_io.m_block_data.data_cnt_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_block_data.data_cnt_q[5] ));
 sky130_fd_sc_hd__nor2_1 \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_X ),
    .Y(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or4_1 \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B  (.A(\m_io.m_block_data.data_cnt_q[2] ),
    .B(\m_io.m_block_data.data_cnt_q[5] ),
    .C(\m_io.m_block_data.data_cnt_q[4] ),
    .D(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_D ),
    .X(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_X ));
 sky130_fd_sc_hd__or4_1 \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_D_sky130_fd_sc_hd__or4_2_X  (.A(\m_io.m_block_data.data_cnt_q[1] ),
    .B(\m_io.m_block_data.data_cnt_q[0] ),
    .C(\m_io.m_block_data.data_cnt_q[3] ),
    .D(net308),
    .X(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__or4_2_B_D ));
 sky130_fd_sc_hd__xor2_1 \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A  (.A(net638),
    .B(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_B ),
    .X(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_io.m_block_data.data_cnt_q[4] ),
    .B(\m_io.m_block_data.data_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor3_2_Y_C ),
    .Y(\m_io.m_block_data.data_cnt_q[5]_sky130_fd_sc_hd__xor2_2_A_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.cfg_cnt_q[0] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_B ),
    .C(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C ),
    .X(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_io.m_config.cfg_cnt_q[0] ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B ),
    .Y(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A ));
 sky130_fd_sc_hd__or2_2 \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B  (.A(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A ),
    .X(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X  (.A(\m_io.m_config.cfg_cnt_q[0] ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C ));
 sky130_fd_sc_hd__and2_1 \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__and2_2_X  (.A(\m_io.m_config.valid_i ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .X(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__nand2_2 \m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A  (.A(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ),
    .Y(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.cfg_cnt_q[1] ));
 sky130_fd_sc_hd__and3b_1 \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X  (.A_N(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_B ),
    .C(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ),
    .X(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N_sky130_fd_sc_hd__and3_2_X  (.A(\m_io.m_config.cfg_cnt_q[1] ),
    .B(\m_io.m_config.cfg_cnt_q[0] ),
    .C(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B ),
    .X(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N ));
 sky130_fd_sc_hd__a31o_1 \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a31o_2_X  (.A1(\m_io.m_config.valid_i ),
    .A2(\m_io.m_config.cfg_cnt_q[0] ),
    .A3(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .B1(\m_io.m_config.cfg_cnt_q[1] ),
    .X(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C ));
 sky130_fd_sc_hd__o311a_1 \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__o311a_2_A1  (.A1(\m_io.m_config.cfg_cnt_q[1] ),
    .A2(\m_io.m_config.cfg_cnt_q[2] ),
    .A3(\m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__nand3_2_C_Y ),
    .B1(\m_io.cmd[2]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .C1(net611),
    .X(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_B ));
 sky130_fd_sc_hd__or3_2 \m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__or3_2_A  (.A(\m_io.m_config.cfg_cnt_q[1] ),
    .B(\m_io.m_config.cfg_cnt_q[2] ),
    .C(\m_io.m_config.cfg_cnt_q[3] ),
    .X(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.cfg_cnt_q[2] ));
 sky130_fd_sc_hd__nor2_1 \m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__and2_1 \m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X  (.A(\m_io.m_config.cfg_cnt_q[2] ),
    .B(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N ),
    .X(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__o21ai_1 \m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y  (.A1(net1852),
    .A2(\m_io.m_config.cfg_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N ),
    .B1(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_B ),
    .Y(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.cfg_cnt_q[3] ));
 sky130_fd_sc_hd__o21a_1 \m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X  (.A1(net1287),
    .A2(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1(\m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__a21boi_1 \m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21boi_2_Y  (.A1(\m_io.m_config.cfg_cnt_q[3] ),
    .A2(\m_io.m_config.cfg_cnt_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B1_N(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_B ),
    .Y(\m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__nand3_1 \m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__nand3_2_C  (.A(\m_io.m_config.valid_i ),
    .B(\m_io.m_config.cfg_cnt_q[0] ),
    .C(\m_io.m_config.cfg_cnt_q[3] ),
    .Y(\m_io.m_config.cfg_cnt_q[3]_sky130_fd_sc_hd__nand3_2_C_Y ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.data_i[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.m_config.data_i[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[0] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net3),
    .X(\m_io.m_config.data_i[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.data_i[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.m_config.data_i[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[1] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(\m_io.en_q ),
    .B(net609),
    .C(net4),
    .X(\m_io.m_config.data_i[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.data_i[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.m_config.data_i[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[2] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net610),
    .C(net5),
    .X(\m_io.m_config.data_i[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.data_i[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.m_config.data_i[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[3] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net610),
    .C(net6),
    .X(\m_io.m_config.data_i[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_4 \m_io.m_config.data_i[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.m_config.data_i[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[4] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net7),
    .X(\m_io.m_config.data_i[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_4 \m_io.m_config.data_i[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_21_clk),
    .D(\m_io.m_config.data_i[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[5] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net8),
    .X(\m_io.m_config.data_i[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_4 \m_io.m_config.data_i[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_22_clk),
    .D(\m_io.m_config.data_i[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[6] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net9),
    .X(\m_io.m_config.data_i[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.data_i[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_config.data_i[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.data_i[7] ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.data_i[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net10),
    .X(\m_io.m_config.data_i[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.kk_q[0] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[0] ),
    .A2(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net612),
    .X(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[8] ),
    .A1(\m_io.m_config.kk_q[0] ),
    .S(net483),
    .X(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.kk_q[0] ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__nor3_1 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y  (.A(\m_io.m_config.cfg_cnt_q[0] ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B ),
    .C(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ),
    .Y(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__nand2_2 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B  (.A(net615),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B ),
    .Y(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_io.m_config.valid_i ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B ));
 sky130_fd_sc_hd__and3_2 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B  (.A(\m_io.m_config.valid_i ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .C(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ),
    .X(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__or3_4 \m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B  (.A(\m_io.m_config.cfg_cnt_q[0] ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B ),
    .C(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ),
    .X(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.kk_q[1] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[1] ),
    .A2(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net612),
    .X(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A  (.A(net1744),
    .Y(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__mux2_1 \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A1(\m_blake2.m_hash256.h_flat[9] ),
    .S(net428),
    .X(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B  (.A(net402),
    .B(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ),
    .Y(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .Y(\m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.kk_q[2] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[2] ),
    .A2(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net611),
    .X(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A  (.A(net1881),
    .Y(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__mux2_1 \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A1(\m_blake2.m_hash256.h_flat[10] ),
    .S(net430),
    .X(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .Y(\m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_11_clk),
    .D(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.kk_q[3] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[3] ),
    .A2(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net612),
    .X(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[11] ),
    .A1(\m_io.m_config.kk_q[3] ),
    .S(net499),
    .X(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B  (.A(net405),
    .B(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X ),
    .Y(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C  (.A(\m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .B(\m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_X ),
    .C(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_B1 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.kk_q[3]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.kk_q[3] ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.kk_q[4] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[4] ),
    .A2(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net614),
    .X(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__mux2_1 \m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1  (.A0(\m_blake2.m_hash256.h_flat[12] ),
    .A1(\m_io.m_config.kk_q[4] ),
    .S(net489),
    .X(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.kk_q[4]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.kk_q[4] ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_10_clk),
    .D(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.kk_q[5] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[5] ),
    .A2(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .B1(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net614),
    .X(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__inv_2 \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A  (.A(\m_io.m_config.kk_q[5] ),
    .Y(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__mux2_1 \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0  (.A0(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y ),
    .A1(\m_blake2.m_hash256.h_flat[13] ),
    .S(net435),
    .X(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A  (.A(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__or3_2_B_X ),
    .Y(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[0] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net890),
    .A2(net163),
    .B1(\m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o2bb2a_1 \m_io.m_config.ll_q[0]_sky130_fd_sc_hd__o2bb2a_2_A1_N  (.A1_N(\m_io.m_config.ll_q[0] ),
    .A2_N(net304),
    .B1(net374),
    .B2(\m_blake2.m_hash256.v_q[12][0] ),
    .X(\m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B2 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[0]_sky130_fd_sc_hd__or2_2_A  (.A(net1025),
    .B(net242),
    .X(\m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(net1779),
    .Q(\m_io.m_config.ll_q[10] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1778),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[10]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[10] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(net1741),
    .Q(\m_io.m_config.ll_q[11] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1740),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[11]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[11] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[12] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net924),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[12]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[12] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_io.m_config.ll_q[13]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[7] ),
    .A2(net262),
    .B1(net306),
    .B2(\m_io.m_config.ll_q[13] ),
    .X(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[13] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net926),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[13]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[13] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[14] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1875),
    .A2(net168),
    .B1(\m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[14]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[14] ),
    .B(net248),
    .X(\m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_io.m_config.ll_q[15]_sky130_fd_sc_hd__a221o_2_B2  (.A1(\m_blake2.m_hash256.v_q[12][15] ),
    .A2(net357),
    .B1(net306),
    .B2(\m_io.m_config.ll_q[15] ),
    .C1(net269),
    .X(\m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[15] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1006),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[15]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[15] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_io.m_config.ll_q[16]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[10] ),
    .A2(net265),
    .B1(net305),
    .B2(\m_io.m_config.ll_q[16] ),
    .X(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[16] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1621),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[16]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[16] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[17] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1122),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[17]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[17] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[18] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1208),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o221a_1 \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[12] ),
    .A2(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ),
    .B1(net240),
    .B2(\m_io.m_config.ll_q[18] ),
    .C1(\m_blake2.m_hash256.v_q[12][18]_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_A2_N ));
 sky130_fd_sc_hd__nand2_2 \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1_sky130_fd_sc_hd__nand2_2_Y  (.A(net463),
    .B(net373),
    .Y(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[18]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[18] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[19] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net878),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[19]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[19] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(net1164),
    .Q(\m_io.m_config.ll_q[1] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1163),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o2bb2a_1 \m_io.m_config.ll_q[1]_sky130_fd_sc_hd__o2bb2a_2_A1_N  (.A1_N(\m_io.m_config.ll_q[1] ),
    .A2_N(net304),
    .B1(net370),
    .B2(\m_blake2.m_hash256.v_q[12][1] ),
    .X(\m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[1]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[1] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_io.m_config.ll_q[20]_sky130_fd_sc_hd__a221o_2_B2  (.A1(\m_blake2.m_hash256.v_q[12][20] ),
    .A2(net352),
    .B1(net307),
    .B2(\m_io.m_config.ll_q[20] ),
    .C1(net269),
    .X(\m_blake2.m_hash256.g_d[20]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[20] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1699),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[20]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[20] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[21] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net938),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[21]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[21] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[22] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net831),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[22]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[22] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[23] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1278),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[23]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[23] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[24] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net942),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[24]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[24] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_io.m_config.ll_q[25]_sky130_fd_sc_hd__a221o_2_B2  (.A1(\m_blake2.m_hash256.v_q[12][25] ),
    .A2(net343),
    .B1(net304),
    .B2(\m_io.m_config.ll_q[25] ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[25] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net994),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[25]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[25] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[25]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_io.m_config.ll_q[26]_sky130_fd_sc_hd__a221o_2_B2  (.A1(\m_blake2.m_hash256.v_q[12][26] ),
    .A2(net348),
    .B1(net304),
    .B2(\m_io.m_config.ll_q[26] ),
    .C1(net268),
    .X(\m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[26] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1069),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[26]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[26] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[27] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1432),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[27]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[27] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[28] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1870),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[28]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[28] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[29] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net873),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[29]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[29] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[2] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net952),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__clkinv_2 \m_io.m_config.ll_q[2]_sky130_fd_sc_hd__inv_2_A  (.A(\m_io.m_config.ll_q[2] ),
    .Y(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__o221a_2_X_B2 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[2]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[2] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[30] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net849),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[30]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[30] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[30]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_io.m_config.ll_q[31]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[25] ),
    .A2(net261),
    .B1(net306),
    .B2(\m_io.m_config.ll_q[31] ),
    .X(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_43_clk),
    .D(\m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[31] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net894),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[31]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[31] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[31]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[32]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[32] ),
    .B(net465),
    .C(net376),
    .X(\m_io.m_config.ll_q[32]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[32] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net941),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[32]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[32] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[33]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[33] ),
    .B(net463),
    .C(net368),
    .X(\m_io.m_config.ll_q[33]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[33] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net881),
    .A2(net163),
    .B1(\m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[33]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[33] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22oi_1 \m_io.m_config.ll_q[34]_sky130_fd_sc_hd__a22oi_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[28] ),
    .A2(net259),
    .B1(net304),
    .B2(\m_io.m_config.ll_q[34] ),
    .Y(\m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__o211a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[34] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net879),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[34]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[34] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22oi_1 \m_io.m_config.ll_q[35]_sky130_fd_sc_hd__a22oi_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[29] ),
    .A2(net264),
    .B1(net307),
    .B2(\m_io.m_config.ll_q[35] ),
    .Y(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__o211a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[35] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1677),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net617),
    .X(\m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[35]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[35] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[36]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[36] ),
    .B(net464),
    .C(net384),
    .X(\m_io.m_config.ll_q[36]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[36] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net853),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[36]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[36] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[37]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[37] ),
    .B(net464),
    .C(net394),
    .X(\m_io.m_config.ll_q[37]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[37] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net995),
    .A2(net168),
    .B1(\m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[37]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[37] ),
    .B(net248),
    .X(\m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[38]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[38] ),
    .B(net464),
    .C(net383),
    .X(\m_io.m_config.ll_q[38]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_46_clk),
    .D(\m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[38] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[46] ),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[38]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[38] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22oi_1 \m_io.m_config.ll_q[39]_sky130_fd_sc_hd__a22oi_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[33] ),
    .A2(net261),
    .B1(net306),
    .B2(\m_io.m_config.ll_q[39] ),
    .Y(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[39] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net855),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[39]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[39] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[39]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_32_clk),
    .D(\m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[3] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1140),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net617),
    .X(\m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__clkinv_2 \m_io.m_config.ll_q[3]_sky130_fd_sc_hd__inv_2_A  (.A(\m_io.m_config.ll_q[3] ),
    .Y(\m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X_B2 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[3]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[3] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[40]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[40] ),
    .B(net465),
    .C(net376),
    .X(\m_io.m_config.ll_q[40]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[40] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1277),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net617),
    .X(\m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[40]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[40] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[40]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[41]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[41] ),
    .B(net463),
    .C(net368),
    .X(\m_io.m_config.ll_q[41]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[41] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net848),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net614),
    .X(\m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[41]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[41] ),
    .B(net243),
    .X(\m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[42]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[42] ),
    .B(\m_blake2.m_hash256.last_block_q ),
    .C(net373),
    .X(\m_io.m_config.ll_q[42]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_26_clk),
    .D(\m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[42] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1240),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net614),
    .X(\m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[42]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[42] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_io.m_config.ll_q[43]_sky130_fd_sc_hd__a221o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[37] ),
    .A2(net265),
    .B1(net305),
    .B2(\m_io.m_config.ll_q[43] ),
    .C1(\m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[43] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1249),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net617),
    .X(\m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[43]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[43] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[44]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[44] ),
    .B(net464),
    .C(net395),
    .X(\m_io.m_config.ll_q[44]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[44] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[52] ),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[44]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[44] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22oi_1 \m_io.m_config.ll_q[45]_sky130_fd_sc_hd__a22oi_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[39] ),
    .A2(net262),
    .B1(net307),
    .B2(\m_io.m_config.ll_q[45] ),
    .Y(\m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(\m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[45] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net839),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[45]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[45] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a211o_1 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_io.m_config.ll_q[46] ),
    .A2(net307),
    .B1(\m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ),
    .C1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ),
    .X(\m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ));
 sky130_fd_sc_hd__nor2_4 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .Y(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__nor3b_4 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__nor3b_2_Y  (.A(net466),
    .B(net469),
    .C_N(net475),
    .Y(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ));
 sky130_fd_sc_hd__or2_2 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A ),
    .B(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ),
    .X(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__and3b_4 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__and3b_2_X  (.A_N(net475),
    .B(net469),
    .C(net466),
    .X(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[46] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net875),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[46]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[46] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[47]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[47] ),
    .B(net464),
    .C(net392),
    .X(\m_io.m_config.ll_q[47]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[47] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net868),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[47]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[47] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22oi_1 \m_io.m_config.ll_q[48]_sky130_fd_sc_hd__a22oi_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[42] ),
    .A2(net265),
    .B1(net305),
    .B2(\m_io.m_config.ll_q[48] ),
    .Y(\m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[48] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[56] ),
    .A2(net164),
    .B1(\m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net617),
    .X(\m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[48]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[48] ),
    .B(net244),
    .X(\m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[49]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[49] ),
    .B(net463),
    .C(net368),
    .X(\m_io.m_config.ll_q[49]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_25_clk),
    .D(\m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[49] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[57] ),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net614),
    .X(\m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[49]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[49] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(net904),
    .Q(\m_io.m_config.ll_q[4] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net903),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o2bb2a_1 \m_io.m_config.ll_q[4]_sky130_fd_sc_hd__o2bb2a_2_A1_N  (.A1_N(\m_io.m_config.ll_q[4] ),
    .A2_N(net307),
    .B1(net384),
    .B2(\m_blake2.m_hash256.v_q[12][4] ),
    .X(\m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[4]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[4] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_io.m_config.ll_q[50]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[44] ),
    .A2(net259),
    .B1(net304),
    .B2(\m_io.m_config.ll_q[50] ),
    .X(\m_io.m_config.ll_q[50]_sky130_fd_sc_hd__a22o_2_B2_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_33_clk),
    .D(\m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[50] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[58] ),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net614),
    .X(\m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[50]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[50] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[51]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[51] ),
    .B(net465),
    .C(net373),
    .X(\m_io.m_config.ll_q[51]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_34_clk),
    .D(\m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[51] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[59] ),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[51]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[51] ),
    .B(net243),
    .X(\m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[52]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[52] ),
    .B(net464),
    .C(net384),
    .X(\m_io.m_config.ll_q[52]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[52] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1146),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[52]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[52] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[52]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[53]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[53] ),
    .B(net464),
    .C(net395),
    .X(\m_io.m_config.ll_q[53]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[53] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net836),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[53]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[53] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[54]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[54] ),
    .B(net464),
    .C(net383),
    .X(\m_io.m_config.ll_q[54]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[54] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net892),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[54]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[54] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[54]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[55]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[55] ),
    .B(net464),
    .C(net392),
    .X(\m_io.m_config.ll_q[55]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[55] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[63] ),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[55]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[55] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a211o_1 \m_io.m_config.ll_q[56]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_io.m_config.ll_q[56] ),
    .A2(net307),
    .B1(\m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ),
    .C1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ),
    .X(\m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_27_clk),
    .D(\m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[56] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[0] ),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net614),
    .X(\m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[56]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[56] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_io.m_config.ll_q[57]_sky130_fd_sc_hd__a221o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[51] ),
    .A2(net259),
    .B1(net304),
    .B2(\m_io.m_config.ll_q[57] ),
    .C1(\m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[57] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[1] ),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net611),
    .X(\m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[57]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[57] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[58]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[58] ),
    .B(net463),
    .C(net373),
    .X(\m_io.m_config.ll_q[58]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[58] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[2] ),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net611),
    .X(\m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[58]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[58] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a221o_1 \m_io.m_config.ll_q[59]_sky130_fd_sc_hd__a221o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[53] ),
    .A2(net260),
    .B1(net305),
    .B2(\m_io.m_config.ll_q[59] ),
    .C1(\m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(\m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A2 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[59] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[3] ),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net611),
    .X(\m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[59]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[59] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_41_clk),
    .D(net912),
    .Q(\m_io.m_config.ll_q[5] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net911),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o2bb2a_1 \m_io.m_config.ll_q[5]_sky130_fd_sc_hd__o2bb2a_2_A1_N  (.A1_N(\m_io.m_config.ll_q[5] ),
    .A2_N(net306),
    .B1(net394),
    .B2(\m_blake2.m_hash256.v_q[12][5] ),
    .X(\m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1 ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[5]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[5] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a211o_1 \m_io.m_config.ll_q[60]_sky130_fd_sc_hd__a211o_2_A1  (.A1(\m_io.m_config.ll_q[60] ),
    .A2(net307),
    .B1(\m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__a2bb2o_2_A1_N_X ),
    .C1(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ),
    .X(\m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_D ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_37_clk),
    .D(\m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[60] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[4] ),
    .A2(net168),
    .B1(\m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net621),
    .X(\m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[60]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[60] ),
    .B(net248),
    .X(\m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[61]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[61] ),
    .B(net465),
    .C(net395),
    .X(\m_io.m_config.ll_q[61]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_38_clk),
    .D(\m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[61] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[5] ),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net621),
    .X(\m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[61]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[61] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.ll_q[62]_sky130_fd_sc_hd__and3_2_A  (.A(\m_io.m_config.ll_q[62] ),
    .B(net464),
    .C(net392),
    .X(\m_io.m_config.ll_q[62]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[62] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[6] ),
    .A2(net166),
    .B1(\m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net619),
    .X(\m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[62]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[62] ),
    .B(net246),
    .X(\m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22oi_1 \m_io.m_config.ll_q[63]_sky130_fd_sc_hd__a22oi_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[57] ),
    .A2(net261),
    .B1(net306),
    .B2(\m_io.m_config.ll_q[63] ),
    .Y(\m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(\m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[63] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[7] ),
    .A2(net162),
    .B1(\m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[63]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[63] ),
    .B(net242),
    .X(\m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_47_clk),
    .D(\m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[6] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net969),
    .A2(net167),
    .B1(\m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net618),
    .X(\m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[6]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[6] ),
    .B(net247),
    .X(\m_io.m_config.ll_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__a22o_1 \m_io.m_config.ll_q[7]_sky130_fd_sc_hd__a22o_2_B2  (.A1(\m_blake2.m_hash256.block_idx_plus_one_q[1] ),
    .A2(net261),
    .B1(net306),
    .B2(\m_io.m_config.ll_q[7] ),
    .X(\m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_42_clk),
    .D(\m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[7] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net1096),
    .A2(net165),
    .B1(\m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net620),
    .X(\m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[7]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[7] ),
    .B(net245),
    .X(\m_io.m_config.ll_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_30_clk),
    .D(net1893),
    .Q(\m_io.m_config.ll_q[8] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.ll_q[16] ),
    .A2(net163),
    .B1(\m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net616),
    .X(\m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[8]_sky130_fd_sc_hd__or2_2_A  (.A(net1892),
    .B(net243),
    .X(\m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_28_clk),
    .D(\m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.ll_q[9] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(net999),
    .A2(net161),
    .B1(\m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net613),
    .X(\m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.ll_q[9]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.ll_q[9] ),
    .B(net241),
    .X(\m_io.m_config.ll_q[9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.nn_q[0] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[0] ),
    .A2(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net611),
    .X(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_2 \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A  (.A(\m_io.m_config.nn_q[0] ),
    .B(net485),
    .Y(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.nn_q[0] ),
    .B(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__nor2_1 \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor2_2_Y  (.A(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_C ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A ),
    .Y(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__or2_2_A_B ));
 sky130_fd_sc_hd__xor2_1 \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A  (.A(\m_io.m_config.nn_q[0] ),
    .B(\m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__xor2_2_B_X ),
    .X(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__or4_1 \m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A  (.A(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A_X ),
    .B(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .C(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .D(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .X(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.nn_q[1] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[1] ),
    .A2(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net612),
    .X(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__inv_2 \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__inv_2_A  (.A(\m_io.m_config.nn_q[1] ),
    .Y(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_io.m_config.nn_q[1] ),
    .B(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_io.m_config.nn_q[1]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_24_clk),
    .D(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.nn_q[2] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[2] ),
    .A2(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net612),
    .X(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__inv_2 \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__inv_2_A  (.A(\m_io.m_config.nn_q[2] ),
    .Y(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_io.m_config.nn_q[2] ),
    .B(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_io.m_config.nn_q[2]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.nn_q[3] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[3] ),
    .A2(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net612),
    .X(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__or2_2_A  (.A(\m_io.m_config.nn_q[3] ),
    .B(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__xnor2_1 \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_io.m_config.nn_q[3] ),
    .B(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ),
    .Y(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ),
    .B(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ),
    .Y(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_blake2.m_hash256.res_cnt_q[3] ),
    .B(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .Y(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_X  (.A(\m_blake2.m_hash256.res_cnt_q[3] ),
    .B(\m_blake2.m_hash256.res_cnt_q[2]_sky130_fd_sc_hd__and2_2_A_X ),
    .X(\m_io.m_config.nn_q[3]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.nn_q[4] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[4] ),
    .A2(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net612),
    .X(\m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__or2_1 \m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__or2_2_X  (.A(\m_io.m_config.nn_q[4] ),
    .B(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(\m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__dfxtp_1 \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_23_clk),
    .D(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.nn_q[5] ));
 sky130_fd_sc_hd__o211a_1 \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X  (.A1(\m_io.m_config.data_i[5] ),
    .A2(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .B1(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ),
    .C1(net611),
    .X(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__nand2_1 \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y  (.A(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y ),
    .B(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_A_sky130_fd_sc_hd__or2_2_B_X ),
    .Y(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1 ));
 sky130_fd_sc_hd__inv_2 \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A  (.A(\m_io.m_config.nn_q[5] ),
    .Y(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__xnor2_1 \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A  (.A(\m_io.m_config.nn_q[5] ),
    .B(\m_blake2.m_hash256.res_cnt_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .Y(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__or4_1 \m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A  (.A(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y ),
    .B(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A_B ),
    .C(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or4_2_A_C ),
    .D(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_X ),
    .X(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__dfxtp_2 \m_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q  (.CLK(clknet_leaf_20_clk),
    .D(\m_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .Q(\m_io.m_config.valid_i ));
 sky130_fd_sc_hd__and3_1 \m_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X  (.A(net1906),
    .B(net609),
    .C(net11),
    .X(\m_io.m_config.valid_i_sky130_fd_sc_hd__dfxtp_2_Q_D ));
 sky130_fd_sc_hd__o21a_1 \m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X  (.A1(\m_blake2.m_hash256.fsm_q[0] ),
    .A2(\m_blake2.m_hash256.fsm_q[3] ),
    .B1(\m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .X(\m_io.ready_v_o ));
 sky130_fd_sc_hd__inv_2 \m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__inv_2_Y  (.A(net606),
    .Y(\m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1 ));
 sky130_fd_sc_hd__mux2_1 \m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__mux2_1_A1  (.A0(net427),
    .A1(\m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1 ),
    .S(\m_blake2.m_hash256.fsm_q[3] ),
    .X(block_last_sky130_fd_sc_hd__a22o_2_B2_A2));
 sky130_fd_sc_hd__conb_1 tt_um_essen_635 (.HI(net635));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_0_clk));
 sky130_fd_sc_hd__conb_1 tt_um_essen_623 (.LO(net623));
 sky130_fd_sc_hd__conb_1 tt_um_essen_624 (.LO(net624));
 sky130_fd_sc_hd__conb_1 tt_um_essen_625 (.LO(net625));
 sky130_fd_sc_hd__conb_1 tt_um_essen_626 (.LO(net626));
 sky130_fd_sc_hd__conb_1 tt_um_essen_627 (.LO(net627));
 sky130_fd_sc_hd__conb_1 tt_um_essen_628 (.LO(net628));
 sky130_fd_sc_hd__buf_2 uio_out_sky130_fd_sc_hd__buf_2_X (.A(\m_io.ready_v_o ),
    .X(uio_out[3]));
 sky130_fd_sc_hd__buf_2 uio_out_sky130_fd_sc_hd__buf_2_X_1 (.A(\m_io.hash_v_o ),
    .X(uio_out[7]));
 sky130_fd_sc_hd__conb_1 tt_um_essen_629 (.LO(net629));
 sky130_fd_sc_hd__conb_1 tt_um_essen_630 (.LO(net630));
 sky130_fd_sc_hd__conb_1 tt_um_essen_631 (.LO(net631));
 sky130_fd_sc_hd__conb_1 tt_um_essen_632 (.LO(net632));
 sky130_fd_sc_hd__conb_1 tt_um_essen_633 (.LO(net633));
 sky130_fd_sc_hd__conb_1 tt_um_essen_634 (.HI(net634));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q (.CLK(clknet_leaf_19_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D),
    .Q(uo_out[7]));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1 (.CLK(clknet_leaf_19_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D),
    .Q(uo_out[6]));
 sky130_fd_sc_hd__a22o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D_sky130_fd_sc_hd__a22o_2_X (.A1(\m_io.m_config.data_i[6] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B2(\hash[6] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2 (.CLK(clknet_leaf_19_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D),
    .Q(uo_out[5]));
 sky130_fd_sc_hd__o22a_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X (.A1(\m_io.m_config.data_i[5] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_B1),
    .B2(\hash[5] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D));
 sky130_fd_sc_hd__clkinv_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__inv_2_Y (.A(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .Y(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_A2));
 sky130_fd_sc_hd__clkinv_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__inv_2_Y (.A(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .Y(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_B1));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3 (.CLK(clknet_leaf_20_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D),
    .Q(uo_out[4]));
 sky130_fd_sc_hd__a22o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D_sky130_fd_sc_hd__a22o_2_X (.A1(\m_io.m_config.data_i[4] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B2(\hash[4] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4 (.CLK(clknet_leaf_19_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D),
    .Q(uo_out[3]));
 sky130_fd_sc_hd__a22o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D_sky130_fd_sc_hd__a22o_2_X (.A1(\m_io.m_config.data_i[3] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B2(\hash[3] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5 (.CLK(clknet_leaf_19_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D),
    .Q(uo_out[2]));
 sky130_fd_sc_hd__a21o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X (.A1(\hash[2] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X_B1),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D));
 sky130_fd_sc_hd__a22o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X (.A1(\m_io.cmd[2] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .B2(\m_io.m_config.data_i[2] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X_B1));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6 (.CLK(clknet_leaf_19_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D),
    .Q(uo_out[1]));
 sky130_fd_sc_hd__a21o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X (.A1(\hash[1] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X_B1),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D));
 sky130_fd_sc_hd__a22o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X (.A1(\m_io.cmd[1] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .B2(\m_io.m_config.data_i[1] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X_B1));
 sky130_fd_sc_hd__dfxtp_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7 (.CLK(clknet_leaf_20_clk),
    .D(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D),
    .Q(uo_out[0]));
 sky130_fd_sc_hd__a21o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X (.A1(\hash[0] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D));
 sky130_fd_sc_hd__a22o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X (.A1(\m_io.m_config.valid_i ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .B2(\m_io.m_config.data_i[0] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1));
 sky130_fd_sc_hd__a22o_1 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X (.A1(\m_io.m_config.data_i[7] ),
    .A2(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .B1(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1),
    .B2(\hash[7] ),
    .X(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D));
 sky130_fd_sc_hd__nor2_2 uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__nor2_2_Y (.A(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2),
    .B(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A2),
    .Y(uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B1));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_2319 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(ena),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(rst_n),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(ui_in[0]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(ui_in[1]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(ui_in[2]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[3]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(ui_in[4]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[5]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[6]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(ui_in[7]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(uio_in[0]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(uio_in[1]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(uio_in[2]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(uio_in[4]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(uio_in[5]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 fanout17 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 fanout19 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__or2_2_A_X ),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 fanout20 (.A(net23),
    .X(net20));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net23),
    .X(net21));
 sky130_fd_sc_hd__buf_4 fanout22 (.A(net23),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(net27),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(net27),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_2 fanout27 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net27));
 sky130_fd_sc_hd__buf_4 fanout28 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_4 fanout30 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 fanout31 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 fanout32 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 fanout33 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 fanout37 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 fanout39 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net39));
 sky130_fd_sc_hd__buf_4 fanout40 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 fanout43 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 fanout47 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 fanout48 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 fanout49 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 fanout51 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 fanout52 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 fanout53 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_4 fanout54 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net54));
 sky130_fd_sc_hd__buf_2 fanout55 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net55));
 sky130_fd_sc_hd__buf_4 fanout56 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 fanout57 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_4 fanout58 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 fanout59 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_4 fanout60 (.A(net63),
    .X(net60));
 sky130_fd_sc_hd__buf_2 fanout61 (.A(net63),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 fanout62 (.A(net63),
    .X(net62));
 sky130_fd_sc_hd__buf_2 fanout63 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_2_Y ),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net64));
 sky130_fd_sc_hd__buf_2 fanout65 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_4 fanout66 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 fanout67 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 fanout69 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_4 fanout70 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 fanout71 (.A(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_4 fanout72 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_2 fanout73 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 fanout75 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 fanout76 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net76));
 sky130_fd_sc_hd__buf_2 fanout77 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 fanout78 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 fanout79 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_4 fanout80 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_2 fanout81 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_4 fanout82 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net82));
 sky130_fd_sc_hd__buf_2 fanout83 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_4 fanout84 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 fanout85 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2_X ),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 fanout89 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2_X ),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_4 fanout90 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2_X ),
    .X(net90));
 sky130_fd_sc_hd__buf_2 fanout91 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_2_X ),
    .X(net91));
 sky130_fd_sc_hd__buf_4 fanout92 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1_X ),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1_X ),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_4 fanout94 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1_X ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_1_X ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 fanout96 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 fanout97 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_2 fanout99 (.A(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net99));
 sky130_fd_sc_hd__buf_6 fanout100 (.A(net103),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(net103),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_2 fanout102 (.A(net103),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__nand4_2_C_Y ),
    .X(net103));
 sky130_fd_sc_hd__buf_4 fanout104 (.A(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_4 fanout105 (.A(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 fanout107 (.A(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_4 fanout108 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ),
    .X(net108));
 sky130_fd_sc_hd__buf_2 fanout109 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_4 fanout110 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 fanout113 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_4 fanout114 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 fanout115 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net116));
 sky130_fd_sc_hd__buf_2 fanout117 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_4 fanout118 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 fanout119 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net123),
    .X(net120));
 sky130_fd_sc_hd__buf_2 fanout121 (.A(net123),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_4 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__buf_2 fanout123 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_X ),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_4 fanout124 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 fanout127 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 fanout129 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4_X ),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4_X ),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 fanout134 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4_X ),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_2 fanout135 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_4_X ),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 fanout136 (.A(net139),
    .X(net136));
 sky130_fd_sc_hd__buf_2 fanout137 (.A(net139),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_4 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_3_X ),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net143),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net143),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_2 fanout143 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_2_X ),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 fanout146 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_2 fanout147 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_4 fanout148 (.A(net151),
    .X(net148));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net151),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_X ),
    .X(net151));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(\m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(net152));
 sky130_fd_sc_hd__buf_4 fanout153 (.A(net154),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 fanout154 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net154));
 sky130_fd_sc_hd__buf_4 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_4 fanout156 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net157));
 sky130_fd_sc_hd__buf_2 fanout158 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 fanout161 (.A(net163),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_2 fanout163 (.A(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net168),
    .X(net164));
 sky130_fd_sc_hd__buf_2 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_2 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__buf_2 fanout168 (.A(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(net168));
 sky130_fd_sc_hd__buf_4 fanout169 (.A(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout170 (.A(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_4 fanout171 (.A(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_8 fanout174 (.A(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ),
    .X(net174));
 sky130_fd_sc_hd__buf_4 fanout175 (.A(\m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B ),
    .X(net175));
 sky130_fd_sc_hd__buf_4 fanout176 (.A(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ),
    .X(net176));
 sky130_fd_sc_hd__buf_4 fanout177 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_4 fanout178 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_4 fanout179 (.A(net180),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_4 fanout180 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ),
    .X(net180));
 sky130_fd_sc_hd__buf_4 fanout181 (.A(net184),
    .X(net181));
 sky130_fd_sc_hd__buf_6 fanout182 (.A(net183),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(net184),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net189),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(net189),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_4 fanout189 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 fanout190 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net190));
 sky130_fd_sc_hd__buf_2 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net193));
 sky130_fd_sc_hd__buf_2 fanout194 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 fanout195 (.A(net197),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_4 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_2 fanout197 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_4 fanout198 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(net200),
    .X(net199));
 sky130_fd_sc_hd__buf_2 fanout200 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(net204),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_4 fanout203 (.A(net204),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_4 fanout204 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_1_Y ),
    .X(net204));
 sky130_fd_sc_hd__buf_4 fanout205 (.A(net208),
    .X(net205));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__buf_4 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__clkbuf_4 fanout208 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(net212),
    .X(net209));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__buf_2 fanout212 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net212));
 sky130_fd_sc_hd__buf_4 fanout213 (.A(net216),
    .X(net213));
 sky130_fd_sc_hd__buf_6 fanout214 (.A(net216),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_1_Y ),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 fanout218 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y ),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_4 fanout222 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(net222));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(net225));
 sky130_fd_sc_hd__buf_2 fanout226 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__buf_4 fanout228 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ),
    .X(net228));
 sky130_fd_sc_hd__buf_4 fanout229 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(net229));
 sky130_fd_sc_hd__buf_2 fanout230 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 fanout231 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 fanout232 (.A(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net234));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 fanout237 (.A(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_4 fanout238 (.A(net239),
    .X(net238));
 sky130_fd_sc_hd__buf_2 fanout239 (.A(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ),
    .X(net239));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ),
    .X(net240));
 sky130_fd_sc_hd__buf_2 fanout241 (.A(net243),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_2 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_2 fanout243 (.A(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 fanout244 (.A(net248),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_2 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(net248),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 fanout248 (.A(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ),
    .X(net248));
 sky130_fd_sc_hd__buf_6 fanout249 (.A(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 fanout250 (.A(net252),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__buf_4 fanout252 (.A(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1_Y ),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(net254),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_8 fanout254 (.A(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ),
    .X(net255));
 sky130_fd_sc_hd__buf_2 fanout256 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_4 fanout260 (.A(net265),
    .X(net260));
 sky130_fd_sc_hd__buf_2 fanout261 (.A(net263),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 fanout262 (.A(net263),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_2 fanout264 (.A(net265),
    .X(net264));
 sky130_fd_sc_hd__buf_2 fanout265 (.A(\m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net265));
 sky130_fd_sc_hd__buf_6 fanout266 (.A(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ),
    .X(net266));
 sky130_fd_sc_hd__buf_6 fanout267 (.A(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2 ),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_4 fanout268 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 fanout269 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_4 fanout273 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net273));
 sky130_fd_sc_hd__buf_6 fanout274 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_8 fanout275 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ),
    .X(net275));
 sky130_fd_sc_hd__buf_2 fanout276 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_4 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_4 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_4 fanout279 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y ),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_4 fanout280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__clkbuf_2 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_2 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y ),
    .X(net283));
 sky130_fd_sc_hd__buf_4 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(net288),
    .X(net287));
 sky130_fd_sc_hd__buf_4 fanout288 (.A(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_4 fanout289 (.A(net290),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_4 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__buf_2 fanout291 (.A(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_4 fanout292 (.A(net294),
    .X(net292));
 sky130_fd_sc_hd__buf_2 fanout293 (.A(net294),
    .X(net293));
 sky130_fd_sc_hd__buf_2 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 fanout295 (.A(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y ),
    .X(net295));
 sky130_fd_sc_hd__buf_4 fanout296 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .X(net296));
 sky130_fd_sc_hd__buf_2 fanout297 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(net299),
    .X(net298));
 sky130_fd_sc_hd__buf_4 fanout299 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ),
    .X(net299));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(net301),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 fanout301 (.A(\m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(net301));
 sky130_fd_sc_hd__buf_4 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__buf_4 fanout303 (.A(\m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X ),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_4 fanout304 (.A(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 fanout305 (.A(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net305));
 sky130_fd_sc_hd__buf_2 fanout306 (.A(net307),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_4 fanout307 (.A(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_4 fanout308 (.A(\m_io.cmd[2]_sky130_fd_sc_hd__o21ai_2_A1_Y ),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_4 fanout309 (.A(net314),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 fanout310 (.A(net314),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_4 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__buf_2 fanout312 (.A(net314),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_4 fanout313 (.A(net314),
    .X(net313));
 sky130_fd_sc_hd__buf_2 fanout314 (.A(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_4 fanout315 (.A(net316),
    .X(net315));
 sky130_fd_sc_hd__buf_2 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__buf_2 fanout317 (.A(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_4 fanout318 (.A(net323),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_4 fanout319 (.A(net320),
    .X(net319));
 sky130_fd_sc_hd__buf_2 fanout320 (.A(net323),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_4 fanout321 (.A(net323),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_4 fanout322 (.A(net323),
    .X(net322));
 sky130_fd_sc_hd__buf_4 fanout323 (.A(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_4 fanout324 (.A(net325),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 fanout325 (.A(net326),
    .X(net325));
 sky130_fd_sc_hd__buf_2 fanout326 (.A(net342),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_4 fanout327 (.A(net330),
    .X(net327));
 sky130_fd_sc_hd__buf_4 fanout328 (.A(net330),
    .X(net328));
 sky130_fd_sc_hd__buf_2 fanout329 (.A(net330),
    .X(net329));
 sky130_fd_sc_hd__buf_2 fanout330 (.A(net342),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_4 fanout331 (.A(net332),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_4 fanout332 (.A(net342),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_4 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 fanout334 (.A(net335),
    .X(net334));
 sky130_fd_sc_hd__buf_4 fanout335 (.A(net342),
    .X(net335));
 sky130_fd_sc_hd__buf_4 fanout336 (.A(net341),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_4 fanout337 (.A(net338),
    .X(net337));
 sky130_fd_sc_hd__buf_2 fanout338 (.A(net341),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_4 fanout339 (.A(net340),
    .X(net339));
 sky130_fd_sc_hd__buf_2 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__buf_2 fanout341 (.A(net342),
    .X(net341));
 sky130_fd_sc_hd__buf_4 fanout342 (.A(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_4 fanout343 (.A(net344),
    .X(net343));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout344 (.A(net345),
    .X(net344));
 sky130_fd_sc_hd__buf_2 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_4 fanout346 (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(net346));
 sky130_fd_sc_hd__buf_2 fanout347 (.A(net349),
    .X(net347));
 sky130_fd_sc_hd__clkbuf_2 fanout348 (.A(net349),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_4 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_4 fanout350 (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(net350));
 sky130_fd_sc_hd__buf_2 fanout351 (.A(net353),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_2 fanout352 (.A(net353),
    .X(net352));
 sky130_fd_sc_hd__buf_2 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_4 fanout354 (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_4 fanout355 (.A(net361),
    .X(net355));
 sky130_fd_sc_hd__buf_2 fanout356 (.A(net361),
    .X(net356));
 sky130_fd_sc_hd__buf_2 fanout357 (.A(net361),
    .X(net357));
 sky130_fd_sc_hd__buf_2 fanout358 (.A(net361),
    .X(net358));
 sky130_fd_sc_hd__buf_2 fanout359 (.A(net361),
    .X(net359));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__buf_2 fanout361 (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ),
    .X(net361));
 sky130_fd_sc_hd__clkbuf_4 fanout362 (.A(net365),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 fanout363 (.A(net365),
    .X(net363));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout364 (.A(net365),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_2 fanout365 (.A(net371),
    .X(net365));
 sky130_fd_sc_hd__buf_2 fanout366 (.A(net371),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_4 fanout367 (.A(net371),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(net369),
    .X(net368));
 sky130_fd_sc_hd__buf_2 fanout369 (.A(net370),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_4 fanout371 (.A(net399),
    .X(net371));
 sky130_fd_sc_hd__buf_2 fanout372 (.A(net399),
    .X(net372));
 sky130_fd_sc_hd__buf_2 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__buf_2 fanout374 (.A(net377),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_2 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_2 fanout377 (.A(net399),
    .X(net377));
 sky130_fd_sc_hd__buf_2 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_4 fanout379 (.A(net385),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_4 fanout380 (.A(net382),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_4 fanout381 (.A(net382),
    .X(net381));
 sky130_fd_sc_hd__buf_2 fanout382 (.A(net385),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net385),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_2 fanout384 (.A(net385),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_4 fanout385 (.A(net399),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_4 fanout386 (.A(net388),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_2 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_4 fanout388 (.A(net391),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_4 fanout389 (.A(net391),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_2 fanout390 (.A(net391),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_2 fanout391 (.A(net398),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(net398),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_2 fanout393 (.A(net398),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_2 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__buf_2 fanout395 (.A(net398),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_4 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_4 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_2 fanout398 (.A(net399),
    .X(net398));
 sky130_fd_sc_hd__buf_4 fanout399 (.A(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__and2b_2_B_X ),
    .X(net399));
 sky130_fd_sc_hd__buf_6 fanout400 (.A(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_4 fanout401 (.A(net403),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_4 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_4 fanout403 (.A(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net403));
 sky130_fd_sc_hd__buf_4 fanout404 (.A(net406),
    .X(net404));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout405 (.A(net406),
    .X(net405));
 sky130_fd_sc_hd__buf_2 fanout406 (.A(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y ),
    .X(net406));
 sky130_fd_sc_hd__buf_6 fanout407 (.A(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A ),
    .X(net407));
 sky130_fd_sc_hd__buf_2 fanout408 (.A(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A ),
    .X(net408));
 sky130_fd_sc_hd__buf_4 fanout409 (.A(net410),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 fanout410 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X ),
    .X(net410));
 sky130_fd_sc_hd__buf_4 fanout411 (.A(net412),
    .X(net411));
 sky130_fd_sc_hd__buf_4 fanout412 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X ),
    .X(net412));
 sky130_fd_sc_hd__buf_4 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__buf_4 fanout414 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X ),
    .X(net414));
 sky130_fd_sc_hd__buf_4 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__buf_4 fanout416 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X ),
    .X(net416));
 sky130_fd_sc_hd__buf_4 fanout417 (.A(net418),
    .X(net417));
 sky130_fd_sc_hd__buf_4 fanout418 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(net418));
 sky130_fd_sc_hd__buf_4 fanout419 (.A(net420),
    .X(net419));
 sky130_fd_sc_hd__buf_4 fanout420 (.A(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X ),
    .X(net420));
 sky130_fd_sc_hd__clkbuf_4 fanout421 (.A(net422),
    .X(net421));
 sky130_fd_sc_hd__buf_2 fanout422 (.A(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ),
    .X(net422));
 sky130_fd_sc_hd__clkbuf_2 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__clkbuf_2 fanout424 (.A(net427),
    .X(net424));
 sky130_fd_sc_hd__clkbuf_2 fanout425 (.A(net427),
    .X(net425));
 sky130_fd_sc_hd__clkbuf_4 fanout426 (.A(net427),
    .X(net426));
 sky130_fd_sc_hd__buf_4 fanout427 (.A(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__nor2_2_B_Y ),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_4 fanout428 (.A(net429),
    .X(net428));
 sky130_fd_sc_hd__buf_2 fanout429 (.A(net431),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_4 fanout430 (.A(net431),
    .X(net430));
 sky130_fd_sc_hd__buf_2 fanout431 (.A(net443),
    .X(net431));
 sky130_fd_sc_hd__buf_2 fanout432 (.A(net434),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_2 fanout433 (.A(net434),
    .X(net433));
 sky130_fd_sc_hd__clkbuf_4 fanout434 (.A(net443),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_4 fanout435 (.A(net443),
    .X(net435));
 sky130_fd_sc_hd__clkbuf_2 fanout436 (.A(net443),
    .X(net436));
 sky130_fd_sc_hd__buf_2 fanout437 (.A(net442),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_2 fanout438 (.A(net442),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_2 fanout439 (.A(net441),
    .X(net439));
 sky130_fd_sc_hd__buf_2 fanout440 (.A(net441),
    .X(net440));
 sky130_fd_sc_hd__clkbuf_4 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_4 fanout442 (.A(net443),
    .X(net442));
 sky130_fd_sc_hd__buf_4 fanout443 (.A(\hash[7]_sky130_fd_sc_hd__and2_2_B_A ),
    .X(net443));
 sky130_fd_sc_hd__buf_2 fanout444 (.A(\m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_A ),
    .X(net444));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout445 (.A(\m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_A ),
    .X(net445));
 sky130_fd_sc_hd__buf_4 fanout446 (.A(net448),
    .X(net446));
 sky130_fd_sc_hd__buf_4 fanout447 (.A(net448),
    .X(net447));
 sky130_fd_sc_hd__clkbuf_8 fanout448 (.A(\m_blake2.m_hash256.shift_hash_q ),
    .X(net448));
 sky130_fd_sc_hd__buf_2 fanout449 (.A(\m_blake2.m_hash256.round_q[9] ),
    .X(net449));
 sky130_fd_sc_hd__clkbuf_2 fanout450 (.A(\m_blake2.m_hash256.round_q[7] ),
    .X(net450));
 sky130_fd_sc_hd__buf_2 fanout451 (.A(net453),
    .X(net451));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 fanout453 (.A(\m_blake2.m_hash256.round_q[6] ),
    .X(net453));
 sky130_fd_sc_hd__buf_2 fanout454 (.A(\m_blake2.m_hash256.round_q[5] ),
    .X(net454));
 sky130_fd_sc_hd__buf_2 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__buf_2 fanout456 (.A(\m_blake2.m_hash256.round_q[4] ),
    .X(net456));
 sky130_fd_sc_hd__buf_2 fanout457 (.A(\m_blake2.m_hash256.round_q[3] ),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_2 fanout458 (.A(\m_blake2.m_hash256.round_q[3] ),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_2 fanout459 (.A(\m_blake2.m_hash256.round_q[2] ),
    .X(net459));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout460 (.A(\m_blake2.m_hash256.round_q[2] ),
    .X(net460));
 sky130_fd_sc_hd__buf_2 fanout461 (.A(\m_blake2.m_hash256.round_q[1] ),
    .X(net461));
 sky130_fd_sc_hd__clkbuf_4 fanout462 (.A(\m_blake2.m_hash256.round_q[0] ),
    .X(net462));
 sky130_fd_sc_hd__clkbuf_4 fanout463 (.A(\m_blake2.m_hash256.last_block_q ),
    .X(net463));
 sky130_fd_sc_hd__buf_2 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__buf_2 fanout465 (.A(\m_blake2.m_hash256.last_block_q ),
    .X(net465));
 sky130_fd_sc_hd__buf_4 fanout466 (.A(\m_blake2.m_hash256.g_idx_q[2] ),
    .X(net466));
 sky130_fd_sc_hd__buf_2 fanout467 (.A(\m_blake2.m_hash256.g_idx_q[2] ),
    .X(net467));
 sky130_fd_sc_hd__buf_2 fanout468 (.A(\m_blake2.m_hash256.g_idx_q[2] ),
    .X(net468));
 sky130_fd_sc_hd__clkbuf_4 fanout469 (.A(net470),
    .X(net469));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_4 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__buf_2 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(\m_blake2.m_hash256.g_idx_q[1] ),
    .X(net473));
 sky130_fd_sc_hd__buf_2 fanout474 (.A(net475),
    .X(net474));
 sky130_fd_sc_hd__buf_4 fanout475 (.A(net476),
    .X(net475));
 sky130_fd_sc_hd__buf_2 fanout476 (.A(net477),
    .X(net476));
 sky130_fd_sc_hd__buf_4 fanout477 (.A(\m_blake2.m_hash256.g_idx_q[0] ),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_4 fanout478 (.A(\m_blake2.m_hash256.fsm_q[4] ),
    .X(net478));
 sky130_fd_sc_hd__clkbuf_2 fanout479 (.A(\m_blake2.m_hash256.fsm_q[4] ),
    .X(net479));
 sky130_fd_sc_hd__buf_4 fanout480 (.A(\m_blake2.m_hash256.fsm_q[4] ),
    .X(net480));
 sky130_fd_sc_hd__clkbuf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__buf_2 fanout482 (.A(\m_blake2.m_hash256.fsm_q[2] ),
    .X(net482));
 sky130_fd_sc_hd__buf_2 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_4 fanout484 (.A(net486),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_4 fanout485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__buf_4 fanout486 (.A(\m_blake2.m_hash256.first_block_q ),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_4 fanout487 (.A(net489),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 fanout488 (.A(net489),
    .X(net488));
 sky130_fd_sc_hd__buf_4 fanout489 (.A(\m_blake2.m_hash256.first_block_q ),
    .X(net489));
 sky130_fd_sc_hd__buf_2 fanout490 (.A(net494),
    .X(net490));
 sky130_fd_sc_hd__buf_2 fanout491 (.A(net493),
    .X(net491));
 sky130_fd_sc_hd__buf_2 fanout492 (.A(net493),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_2 fanout493 (.A(net494),
    .X(net493));
 sky130_fd_sc_hd__clkbuf_4 fanout494 (.A(\m_blake2.m_hash256.first_block_q ),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_4 fanout495 (.A(net497),
    .X(net495));
 sky130_fd_sc_hd__buf_2 fanout496 (.A(net497),
    .X(net496));
 sky130_fd_sc_hd__clkbuf_2 fanout497 (.A(net500),
    .X(net497));
 sky130_fd_sc_hd__buf_2 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_4 fanout499 (.A(net500),
    .X(net499));
 sky130_fd_sc_hd__buf_2 fanout500 (.A(\m_blake2.m_hash256.first_block_q ),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_4 fanout501 (.A(net502),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_2 fanout502 (.A(net509),
    .X(net502));
 sky130_fd_sc_hd__clkbuf_4 fanout503 (.A(net504),
    .X(net503));
 sky130_fd_sc_hd__buf_2 fanout504 (.A(net509),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_4 fanout505 (.A(net509),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_4 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__buf_2 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_4 fanout508 (.A(net509),
    .X(net508));
 sky130_fd_sc_hd__buf_2 fanout509 (.A(net539),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_4 fanout510 (.A(net511),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_4 fanout511 (.A(net539),
    .X(net511));
 sky130_fd_sc_hd__clkbuf_4 fanout512 (.A(net516),
    .X(net512));
 sky130_fd_sc_hd__buf_2 fanout513 (.A(net516),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_4 fanout514 (.A(net515),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_4 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_2 fanout516 (.A(net539),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_4 fanout517 (.A(net519),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_2 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__buf_2 fanout519 (.A(net524),
    .X(net519));
 sky130_fd_sc_hd__clkbuf_4 fanout520 (.A(net524),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_2 fanout521 (.A(net524),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_4 fanout522 (.A(net524),
    .X(net522));
 sky130_fd_sc_hd__buf_2 fanout523 (.A(net524),
    .X(net523));
 sky130_fd_sc_hd__buf_2 fanout524 (.A(net539),
    .X(net524));
 sky130_fd_sc_hd__clkbuf_4 fanout525 (.A(net526),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_4 fanout526 (.A(net538),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_4 fanout527 (.A(net529),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_2 fanout528 (.A(net529),
    .X(net528));
 sky130_fd_sc_hd__buf_2 fanout529 (.A(net530),
    .X(net529));
 sky130_fd_sc_hd__clkbuf_4 fanout530 (.A(net538),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_4 fanout531 (.A(net538),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_2 fanout532 (.A(net538),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_4 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__buf_2 fanout534 (.A(net537),
    .X(net534));
 sky130_fd_sc_hd__clkbuf_4 fanout535 (.A(net537),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_2 fanout536 (.A(net537),
    .X(net536));
 sky130_fd_sc_hd__clkbuf_2 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__clkbuf_4 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__buf_4 fanout539 (.A(\m_blake2.m_hash256.f_finished_q ),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(net542),
    .X(net540));
 sky130_fd_sc_hd__clkbuf_2 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_4 fanout542 (.A(net546),
    .X(net542));
 sky130_fd_sc_hd__clkbuf_4 fanout543 (.A(net545),
    .X(net543));
 sky130_fd_sc_hd__clkbuf_2 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__clkbuf_4 fanout545 (.A(net546),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_2 fanout546 (.A(net608),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(net548),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_4 fanout548 (.A(net550),
    .X(net548));
 sky130_fd_sc_hd__clkbuf_4 fanout549 (.A(net550),
    .X(net549));
 sky130_fd_sc_hd__buf_2 fanout550 (.A(net608),
    .X(net550));
 sky130_fd_sc_hd__clkbuf_4 fanout551 (.A(net553),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_2 fanout552 (.A(net553),
    .X(net552));
 sky130_fd_sc_hd__buf_2 fanout553 (.A(net561),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_4 fanout554 (.A(net555),
    .X(net554));
 sky130_fd_sc_hd__clkbuf_4 fanout555 (.A(net561),
    .X(net555));
 sky130_fd_sc_hd__clkbuf_2 fanout556 (.A(net561),
    .X(net556));
 sky130_fd_sc_hd__clkbuf_4 fanout557 (.A(net561),
    .X(net557));
 sky130_fd_sc_hd__buf_2 fanout558 (.A(net561),
    .X(net558));
 sky130_fd_sc_hd__clkbuf_4 fanout559 (.A(net560),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_4 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__clkbuf_2 fanout561 (.A(net608),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_4 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_4 fanout563 (.A(net564),
    .X(net563));
 sky130_fd_sc_hd__buf_2 fanout564 (.A(net567),
    .X(net564));
 sky130_fd_sc_hd__clkbuf_4 fanout565 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_4 fanout566 (.A(net567),
    .X(net566));
 sky130_fd_sc_hd__clkbuf_2 fanout567 (.A(net579),
    .X(net567));
 sky130_fd_sc_hd__clkbuf_4 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(net570),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_2 fanout570 (.A(net571),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_4 fanout571 (.A(net579),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_4 fanout572 (.A(net575),
    .X(net572));
 sky130_fd_sc_hd__clkbuf_4 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_4 fanout574 (.A(net575),
    .X(net574));
 sky130_fd_sc_hd__clkbuf_2 fanout575 (.A(net579),
    .X(net575));
 sky130_fd_sc_hd__clkbuf_4 fanout576 (.A(net578),
    .X(net576));
 sky130_fd_sc_hd__buf_2 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__clkbuf_4 fanout578 (.A(net579),
    .X(net578));
 sky130_fd_sc_hd__buf_2 fanout579 (.A(net608),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_4 fanout580 (.A(net582),
    .X(net580));
 sky130_fd_sc_hd__clkbuf_2 fanout581 (.A(net582),
    .X(net581));
 sky130_fd_sc_hd__clkbuf_2 fanout582 (.A(net590),
    .X(net582));
 sky130_fd_sc_hd__clkbuf_4 fanout583 (.A(net585),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_2 fanout584 (.A(net585),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_4 fanout585 (.A(net590),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_4 fanout586 (.A(net589),
    .X(net586));
 sky130_fd_sc_hd__clkbuf_4 fanout587 (.A(net589),
    .X(net587));
 sky130_fd_sc_hd__clkbuf_4 fanout588 (.A(net589),
    .X(net588));
 sky130_fd_sc_hd__clkbuf_2 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_2 fanout590 (.A(net608),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_4 fanout591 (.A(net592),
    .X(net591));
 sky130_fd_sc_hd__buf_2 fanout592 (.A(net594),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_4 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_2 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__clkbuf_4 fanout595 (.A(net599),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_4 fanout596 (.A(net599),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_2 fanout597 (.A(net599),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_4 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout599 (.A(net608),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_4 fanout600 (.A(net602),
    .X(net600));
 sky130_fd_sc_hd__clkbuf_4 fanout601 (.A(net602),
    .X(net601));
 sky130_fd_sc_hd__buf_2 fanout602 (.A(net603),
    .X(net602));
 sky130_fd_sc_hd__clkbuf_4 fanout603 (.A(net607),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_4 fanout604 (.A(net605),
    .X(net604));
 sky130_fd_sc_hd__clkbuf_4 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__clkbuf_4 fanout606 (.A(net607),
    .X(net606));
 sky130_fd_sc_hd__clkbuf_2 fanout607 (.A(net608),
    .X(net607));
 sky130_fd_sc_hd__buf_2 fanout608 (.A(data_v),
    .X(net608));
 sky130_fd_sc_hd__clkbuf_2 fanout609 (.A(net610),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_2 fanout610 (.A(net615),
    .X(net610));
 sky130_fd_sc_hd__buf_2 fanout611 (.A(net612),
    .X(net611));
 sky130_fd_sc_hd__buf_2 fanout612 (.A(net615),
    .X(net612));
 sky130_fd_sc_hd__buf_2 fanout613 (.A(net614),
    .X(net613));
 sky130_fd_sc_hd__buf_2 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__clkbuf_2 fanout615 (.A(net2),
    .X(net615));
 sky130_fd_sc_hd__buf_2 fanout616 (.A(net621),
    .X(net616));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout617 (.A(net621),
    .X(net617));
 sky130_fd_sc_hd__buf_2 fanout618 (.A(net621),
    .X(net618));
 sky130_fd_sc_hd__buf_2 fanout619 (.A(net620),
    .X(net619));
 sky130_fd_sc_hd__buf_2 fanout620 (.A(net621),
    .X(net620));
 sky130_fd_sc_hd__buf_2 fanout621 (.A(net2),
    .X(net621));
 sky130_fd_sc_hd__conb_1 tt_um_essen_622 (.LO(net622));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_1_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_3_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_4_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_5_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_6_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_7_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_8_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_9_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_10_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_12_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_13_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_15_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_16_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_18_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_19_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_20_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_20_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_21_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_21_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_22_clk (.A(clknet_3_2_0_clk),
    .X(clknet_leaf_22_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_23_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_23_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_24_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_24_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_25_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_25_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_26_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_26_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_27_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_27_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_28_clk (.A(clknet_3_3_0_clk),
    .X(clknet_leaf_28_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_29_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_29_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_30_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_30_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_31_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_31_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_32_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_33_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_33_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_34_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_34_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_35_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_35_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_36_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_36_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_37_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_37_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_38_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_38_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_39_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_39_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_40_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_40_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_41_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_41_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_42_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_42_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_43_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_43_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_44_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_44_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_45_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_45_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_46_clk (.A(clknet_3_7_0_clk),
    .X(clknet_leaf_46_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_47_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_47_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_48_clk (.A(clknet_3_6_0_clk),
    .X(clknet_leaf_48_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_49_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_49_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_50_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_50_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_51_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_51_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_52_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_52_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_53_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_53_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_54_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_55_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_56_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_56_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_57_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_57_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_58_clk (.A(clknet_3_5_0_clk),
    .X(clknet_leaf_58_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_59_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_59_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_60_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_60_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_61_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_61_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_62_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_62_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_63_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_63_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_64_clk (.A(clknet_3_4_0_clk),
    .X(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_65_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_66_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_66_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_67_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_68_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_68_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_69_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_69_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_70_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_70_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_71_clk (.A(clknet_3_1_0_clk),
    .X(clknet_leaf_71_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_72_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_72_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_73_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_73_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_74_clk (.A(clknet_3_0_0_clk),
    .X(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_clk (.A(clknet_0_clk),
    .X(clknet_3_0_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_clk (.A(clknet_0_clk),
    .X(clknet_3_1_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_clk (.A(clknet_0_clk),
    .X(clknet_3_2_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_clk (.A(clknet_0_clk),
    .X(clknet_3_3_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_clk (.A(clknet_0_clk),
    .X(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_clk (.A(clknet_0_clk),
    .X(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_clk (.A(clknet_0_clk),
    .X(clknet_3_6_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_clk (.A(clknet_0_clk),
    .X(clknet_3_7_0_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_3_1_0_clk));
 sky130_fd_sc_hd__inv_6 clkload1 (.A(clknet_3_3_0_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_3_4_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload3 (.A(clknet_3_5_0_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload4 (.A(clknet_3_6_0_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_3_7_0_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload6 (.A(clknet_leaf_2_clk));
 sky130_fd_sc_hd__clkinv_2 clkload7 (.A(clknet_leaf_5_clk));
 sky130_fd_sc_hd__bufinv_16 clkload8 (.A(clknet_leaf_7_clk));
 sky130_fd_sc_hd__inv_8 clkload9 (.A(clknet_leaf_74_clk));
 sky130_fd_sc_hd__clkinv_8 clkload10 (.A(clknet_leaf_65_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload11 (.A(clknet_leaf_67_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload12 (.A(clknet_leaf_70_clk));
 sky130_fd_sc_hd__inv_6 clkload13 (.A(clknet_leaf_14_clk));
 sky130_fd_sc_hd__clkinv_2 clkload14 (.A(clknet_leaf_17_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload15 (.A(clknet_leaf_21_clk));
 sky130_fd_sc_hd__inv_6 clkload16 (.A(clknet_leaf_22_clk));
 sky130_fd_sc_hd__inv_8 clkload17 (.A(clknet_leaf_11_clk));
 sky130_fd_sc_hd__clkbuf_8 clkload18 (.A(clknet_leaf_24_clk));
 sky130_fd_sc_hd__inv_8 clkload19 (.A(clknet_leaf_27_clk));
 sky130_fd_sc_hd__inv_12 clkload20 (.A(clknet_leaf_49_clk));
 sky130_fd_sc_hd__inv_16 clkload21 (.A(clknet_leaf_50_clk));
 sky130_fd_sc_hd__inv_4 clkload22 (.A(clknet_leaf_62_clk));
 sky130_fd_sc_hd__inv_16 clkload23 (.A(clknet_leaf_63_clk));
 sky130_fd_sc_hd__inv_16 clkload24 (.A(clknet_leaf_64_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload25 (.A(clknet_leaf_45_clk));
 sky130_fd_sc_hd__inv_8 clkload26 (.A(clknet_leaf_51_clk));
 sky130_fd_sc_hd__inv_12 clkload27 (.A(clknet_leaf_54_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload28 (.A(clknet_leaf_55_clk));
 sky130_fd_sc_hd__clkinv_2 clkload29 (.A(clknet_leaf_29_clk));
 sky130_fd_sc_hd__inv_8 clkload30 (.A(clknet_leaf_31_clk));
 sky130_fd_sc_hd__inv_8 clkload31 (.A(clknet_leaf_32_clk));
 sky130_fd_sc_hd__clkinv_2 clkload32 (.A(clknet_leaf_35_clk));
 sky130_fd_sc_hd__inv_8 clkload33 (.A(clknet_leaf_36_clk));
 sky130_fd_sc_hd__inv_6 clkload34 (.A(clknet_leaf_46_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\m_io.m_block_data.data_cnt_q[1] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\m_io.m_block_data.data_cnt_q[3] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\m_io.m_block_data.data_cnt_q[5] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\m_io.m_block_data.data_cnt_q[4] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\m_io.m_block_data.data_cnt_q[0] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\m_io.m_block_data.data_cnt_q[2] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\data[3] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\m_blake2.m_hash256.m_matrix[15][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\data[0] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\m_blake2.m_hash256.h_flat[255] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\m_blake2.m_hash256.m_matrix[15][24] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\data[1] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(block_first),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\m_blake2.m_hash256.m_matrix[15][25] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\data[2] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\m_blake2.m_hash256.m_matrix[15][26] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\m_blake2.m_hash256.h_flat[197] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\m_blake2.m_hash256.h_flat[199] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\m_blake2.m_hash256.h_flat[162] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(block_last),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\m_blake2.m_hash256.fsm_q[1] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\m_blake2.m_hash256.h_flat[174] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\m_blake2.m_hash256.h_flat[167] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\m_blake2.m_hash256.h_flat[219] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\m_blake2.m_hash256.h_flat[82] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\m_blake2.m_hash256.h_flat[148] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\m_blake2.m_hash256.h_flat[151] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\m_blake2.m_hash256.h_flat[55] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\m_blake2.m_hash256.h_flat[184] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\m_blake2.m_hash256.h_flat[143] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\m_blake2.m_hash256.h_flat[173] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\m_blake2.m_hash256.h_flat[145] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\m_blake2.m_hash256.h_flat[216] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\m_blake2.m_hash256.h_flat[251] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\m_blake2.m_hash256.h_flat[71] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\m_blake2.m_hash256.h_flat[154] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\m_blake2.m_hash256.h_flat[35] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\m_blake2.m_hash256.h_flat[40] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\m_blake2.m_hash256.h_flat[46] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\m_blake2.m_hash256.h_flat[190] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\m_blake2.m_hash256.h_flat[67] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\m_blake2.m_hash256.h_flat[202] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\m_blake2.m_hash256.h_flat[51] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\m_blake2.m_hash256.h_flat[119] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\m_blake2.m_hash256.h_flat[227] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\m_blake2.m_hash256.h_flat[87] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\m_blake2.m_hash256.h_flat[191] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\m_blake2.m_hash256.h_flat[31] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\m_blake2.m_hash256.h_flat[126] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\m_blake2.m_hash256.h_flat[62] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\m_blake2.m_hash256.h_flat[33] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\m_blake2.m_hash256.h_flat[27] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\m_blake2.m_hash256.h_flat[164] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\m_blake2.m_hash256.h_flat[74] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\m_blake2.m_hash256.h_flat[36] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\m_blake2.m_hash256.h_flat[123] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\m_blake2.m_hash256.h_flat[207] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\m_blake2.m_hash256.h_flat[237] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\m_blake2.m_hash256.h_flat[22] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\m_blake2.m_hash256.h_flat[99] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\m_blake2.m_hash256.h_flat[103] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\m_blake2.m_hash256.h_flat[218] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\m_blake2.m_hash256.h_flat[156] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\m_blake2.m_hash256.h_flat[205] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\m_blake2.m_hash256.h_flat[146] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\m_blake2.m_hash256.h_flat[240] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\m_blake2.m_hash256.h_flat[54] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\m_blake2.m_hash256.h_flat[9] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\m_blake2.m_hash256.h_flat[106] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\m_blake2.m_hash256.h_flat[152] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\m_blake2.m_hash256.h_flat[94] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\m_blake2.m_hash256.h_flat[37] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\m_blake2.m_hash256.h_flat[226] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\m_blake2.m_hash256.h_flat[95] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\m_blake2.m_hash256.h_flat[81] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\m_blake2.m_hash256.h_flat[193] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\m_blake2.m_hash256.h_flat[10] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\m_blake2.m_hash256.h_flat[14] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\m_blake2.m_hash256.h_flat[115] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\m_blake2.m_hash256.h_flat[97] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\m_blake2.m_hash256.h_flat[223] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\m_blake2.m_hash256.h_flat[158] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\m_blake2.m_hash256.h_flat[23] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\m_blake2.m_hash256.h_flat[157] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\m_blake2.m_hash256.h_flat[38] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\m_blake2.m_hash256.h_flat[153] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\m_blake2.m_hash256.h_flat[233] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\m_blake2.m_hash256.h_flat[39] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\m_blake2.m_hash256.h_flat[77] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\m_blake2.m_hash256.h_flat[149] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\m_blake2.m_hash256.h_flat[178] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\m_blake2.m_hash256.h_flat[18] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\m_blake2.m_hash256.h_flat[107] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\m_blake2.m_hash256.h_flat[165] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\m_blake2.m_hash256.h_flat[170] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\m_blake2.m_hash256.h_flat[8] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\m_blake2.m_hash256.h_flat[249] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\m_blake2.m_hash256.h_flat[59] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\m_blake2.m_hash256.h_flat[100] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\m_blake2.m_hash256.h_flat[155] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\m_blake2.m_hash256.h_flat[177] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\m_blake2.m_hash256.h_flat[169] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\m_blake2.m_hash256.h_flat[196] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\m_blake2.m_hash256.h_flat[110] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\m_blake2.m_hash256.h_flat[163] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\m_blake2.m_hash256.h_flat[114] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\m_blake2.m_hash256.h_flat[138] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\m_blake2.m_hash256.h_flat[91] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\m_blake2.m_hash256.h_flat[104] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\m_blake2.m_hash256.h_flat[45] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\m_blake2.m_hash256.h_flat[69] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\m_blake2.m_hash256.h_flat[217] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\m_blake2.m_hash256.h_flat[239] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\m_blake2.m_hash256.h_flat[58] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\m_blake2.m_hash256.h_flat[98] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\m_blake2.m_hash256.h_flat[117] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\m_blake2.m_hash256.h_flat[209] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\m_blake2.m_hash256.h_flat[241] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\m_blake2.m_hash256.h_flat[238] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\m_blake2.m_hash256.h_flat[85] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\m_blake2.m_hash256.h_flat[234] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\m_blake2.m_hash256.h_flat[72] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\m_blake2.m_hash256.h_flat[248] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\m_blake2.m_hash256.h_flat[181] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\m_blake2.m_hash256.h_flat[215] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\m_blake2.m_hash256.h_flat[116] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\m_blake2.m_hash256.h_flat[140] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\m_blake2.m_hash256.h_flat[176] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\m_blake2.m_hash256.h_flat[213] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\m_blake2.m_hash256.h_flat[12] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\m_blake2.m_hash256.h_flat[210] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\m_blake2.m_hash256.h_flat[137] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\m_blake2.m_hash256.h_flat[26] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\m_blake2.m_hash256.m_matrix[0][0] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\m_blake2.m_hash256.h_flat[185] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\m_blake2.m_hash256.h_flat[52] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\m_blake2.m_hash256.h_flat[65] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\m_blake2.m_hash256.h_flat[49] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\m_blake2.m_hash256.h_flat[254] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\m_blake2.m_hash256.h_flat[34] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\m_blake2.m_hash256.h_flat[102] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\m_blake2.m_hash256.h_flat[236] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\m_blake2.m_hash256.h_flat[11] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\m_blake2.m_hash256.h_flat[53] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\m_blake2.m_hash256.h_flat[171] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\m_blake2.m_hash256.h_flat[78] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\m_blake2.m_hash256.h_flat[16] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\m_blake2.m_hash256.h_flat[68] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\m_blake2.m_hash256.h_flat[200] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\m_blake2.m_hash256.h_flat[141] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\m_blake2.m_hash256.h_flat[187] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\m_blake2.m_hash256.h_flat[61] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\m_blake2.m_hash256.h_flat[231] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\m_blake2.m_hash256.h_flat[84] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\m_blake2.m_hash256.h_flat[83] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\m_blake2.m_hash256.h_flat[168] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\m_blake2.m_hash256.h_flat[101] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\m_blake2.m_hash256.h_flat[90] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[57] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\m_blake2.m_hash256.h_flat[20] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\m_blake2.m_hash256.m_matrix[0][6] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\m_blake2.m_hash256.h_flat[201] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\m_blake2.m_hash256.h_flat[203] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\m_blake2.m_hash256.h_flat[111] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\m_blake2.m_hash256.h_flat[147] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\m_blake2.m_hash256.h_flat[60] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\m_blake2.m_hash256.h_flat[228] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\m_blake2.m_hash256.h_flat[189] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\m_blake2.m_hash256.h_flat[142] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\m_blake2.m_hash256.h_flat[21] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\m_blake2.m_hash256.h_flat[235] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\m_blake2.m_hash256.h_flat[161] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\m_blake2.m_hash256.h_flat[225] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\m_blake2.m_hash256.h_flat[247] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\m_blake2.m_hash256.h_flat[66] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\m_blake2.m_hash256.h_flat[42] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\data[4] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\m_blake2.m_hash256.h_flat[113] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\m_blake2.m_hash256.h_flat[175] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\m_blake2.m_hash256.h_flat[80] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\m_blake2.m_hash256.h_flat[63] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\m_blake2.m_hash256.h_flat[118] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\m_blake2.m_hash256.fsm_q[0] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\m_blake2.m_hash256.slow_output_q_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\m_blake2.m_hash256.h_flat[43] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\m_blake2.m_hash256.h_flat[127] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\m_blake2.m_hash256.v_q[15][30] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\m_blake2.m_hash256.h_flat[41] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\m_blake2.m_hash256.h_flat[206] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\m_blake2.m_hash256.h_flat[186] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\m_blake2.m_hash256.m_matrix[1][18] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\m_blake2.m_hash256.m_matrix[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\m_blake2.m_hash256.h_flat[86] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\m_io.m_config.ll_q[30] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\m_blake2.m_hash256.h_flat[47] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\m_blake2.m_hash256.h_flat[109] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\data[6] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\m_blake2.m_hash256.h_flat[30] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\m_io.m_config.ll_q[61] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\m_blake2.m_hash256.h_flat[139] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\m_blake2.m_hash256.h_flat[245] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\m_io.m_config.ll_q[53] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\m_blake2.m_hash256.h_flat[75] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\m_blake2.m_hash256.h_flat[221] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\m_blake2.m_hash256.h_flat[13] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\m_blake2.m_hash256.h_flat[136] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\m_blake2.m_hash256.v_q[4][9] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\m_blake2.m_hash256.h_flat[17] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\m_blake2.m_hash256.h_flat[222] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\m_blake2.m_hash256.h_flat[122] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\m_io.m_config.ll_q[49] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\m_io.m_config.ll_q[38] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\m_blake2.m_hash256.h_flat[195] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\m_blake2.m_hash256.slow_output_q ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\m_io.m_config.ll_q[44] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\m_blake2.m_hash256.h_flat[70] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\m_io.m_config.ll_q[47] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\m_blake2.m_hash256.v_q[4][13] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\m_blake2.m_hash256.h_flat[96] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\m_blake2.m_hash256.v_q[15][10] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\m_blake2.m_hash256.h_flat[242] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\m_blake2.m_hash256.h_flat[121] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\m_blake2.m_hash256.v_q[14][16] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\m_blake2.m_hash256.h_flat[79] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\m_blake2.m_hash256.h_flat[182] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\m_blake2.m_hash256.h_flat[57] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\m_blake2.m_hash256.h_flat[183] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\m_blake2.m_hash256.h_flat[15] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\m_blake2.m_hash256.v_q[4][30] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\m_io.m_config.ll_q[55] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\m_blake2.m_hash256.v_q[4][7] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\m_blake2.m_hash256.m_matrix[0][3] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\m_blake2.m_hash256.h_flat[135] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\m_io.m_config.ll_q[37] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\data[7] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\m_io.m_config.ll_q[54] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\m_blake2.m_hash256.v_q[10][21] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\m_blake2.m_hash256.v_q[5][11] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\m_io.m_config.ll_q[27] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\m_io.m_config.ll_q[42] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\m_blake2.m_hash256.v_q[4][27] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\m_io.m_config.ll_q[41] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\m_blake2.m_hash256.v_q[15][8] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\m_blake2.m_hash256.v_q[4][18] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\m_blake2.m_hash256.h_flat[89] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\m_blake2.m_hash256.h_flat[232] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\m_blake2.m_hash256.v_q[4][19] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\m_blake2.m_hash256.h_flat[108] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\m_blake2.m_hash256.h_flat[92] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\m_blake2.m_hash256.v_q[4][26] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\m_io.m_config.ll_q[8] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\m_blake2.m_hash256.v_q[4][21] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\m_io.m_config.ll_q[62] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\m_blake2.m_hash256.h_flat[48] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\m_io.m_config.ll_q[39] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\m_blake2.m_hash256.v_q[1][11] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\m_blake2.m_hash256.h_flat[93] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\m_blake2.m_hash256.v_q[9][24] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\m_blake2.m_hash256.v_q[15][22] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\m_blake2.m_hash256.h_flat[180] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\m_blake2.m_hash256.h_flat[244] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\m_blake2.m_hash256.v_q[4][17] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\m_blake2.m_hash256.v_q[4][23] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\m_io.m_config.ll_q[12] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\m_io.m_config.ll_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\m_blake2.m_hash256.v_q[6][1] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\m_blake2.m_hash256.v_q[4][11] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\m_blake2.m_hash256.v_q[4][15] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\m_blake2.m_hash256.h_flat[192] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\m_blake2.m_hash256.h_flat[73] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\m_blake2.m_hash256.v_q[14][20] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\m_io.m_config.ll_q[13] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\m_io.m_config.ll_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\m_blake2.m_hash256.h_flat[229] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\m_blake2.m_hash256.v_q[0][17] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\m_blake2.m_hash256.h_flat[76] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\m_blake2.m_hash256.v_q[10][1] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\m_blake2.m_hash256.v_q[2][11] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\m_blake2.m_hash256.v_q[4][25] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\m_blake2.m_hash256.v_q[4][31] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\m_blake2.m_hash256.v_q[13][24] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\m_blake2.m_hash256.v_q[6][3] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\m_blake2.m_hash256.v_q[1][17] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\m_blake2.m_hash256.h_flat[50] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\m_io.m_config.ll_q[20] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\m_blake2.m_hash256.h_flat[105] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\m_io.m_config.ll_q[21] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\m_blake2.m_hash256.v_q[9][20] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\m_blake2.m_hash256.v_q[4][10] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\m_blake2.m_hash256.v_q[4][29] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\m_blake2.m_hash256.v_q[4][14] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\m_blake2.m_hash256.v_q[6][21] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\m_blake2.m_hash256.v_q[5][25] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\m_blake2.m_hash256.v_q[6][22] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\m_blake2.m_hash256.v_q[4][16] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\m_blake2.m_hash256.m_matrix[15][31] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\m_blake2.m_hash256.v_q[4][20] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\m_blake2.m_hash256.v_q[5][31] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\m_io.m_config.ll_q[29] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\m_blake2.m_hash256.v_q[6][18] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\m_blake2.m_hash256.v_q[9][28] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\m_io.m_config.ll_q[40] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\m_io.m_config.ll_q[32] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\m_blake2.m_hash256.v_q[14][27] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\m_blake2.m_hash256.v_q[6][30] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\m_blake2.m_hash256.v_q[6][5] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\m_blake2.m_hash256.m_matrix[0][2] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\m_blake2.m_hash256.v_q[6][0] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\m_blake2.m_hash256.v_q[0][28] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\m_blake2.m_hash256.v_q[0][5] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\m_blake2.m_hash256.v_q[6][4] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\m_io.m_config.ll_q[10] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\m_blake2.m_hash256.v_q[3][11] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\m_blake2.m_hash256.m_matrix[12][10] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\m_blake2.m_hash256.v_q[6][27] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\m_blake2.m_hash256.v_q[3][18] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\m_blake2.m_hash256.v_q[6][10] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\m_blake2.m_hash256.v_q[10][28] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\m_blake2.m_hash256.v_q[4][22] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\m_blake2.m_hash256.v_q[0][20] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\m_blake2.m_hash256.v_q[4][8] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\m_blake2.m_hash256.v_q[3][17] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\m_blake2.m_hash256.m_matrix[5][13] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\m_blake2.m_hash256.h_flat[212] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\m_blake2.m_hash256.v_q[1][0] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\m_blake2.m_hash256.m_matrix[10][3] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\m_blake2.m_hash256.v_q[0][27] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\m_blake2.m_hash256.v_q[3][10] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\m_io.m_config.ll_q[14] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\m_blake2.m_hash256.v_q[0][18] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\m_blake2.m_hash256.v_q[5][4] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\m_blake2.m_hash256.v_q[5][5] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\m_blake2.m_hash256.v_q[0][26] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\m_blake2.m_hash256.v_q[0][6] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\m_blake2.m_hash256.v_q[3][9] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\m_blake2.m_hash256.v_q[3][24] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\m_blake2.m_hash256.v_q[5][28] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\m_blake2.m_hash256.v_q[5][2] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\m_blake2.m_hash256.v_q[1][2] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\m_blake2.m_hash256.v_q[0][16] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\m_blake2.m_hash256.m_matrix[6][30] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\m_blake2.m_hash256.v_q[6][26] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\m_blake2.m_hash256.v_q[12][4] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\m_blake2.m_hash256.v_q[0][3] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\m_blake2.m_hash256.v_q[4][6] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\m_blake2.m_hash256.m_matrix[0][25] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\m_blake2.m_hash256.v_q[6][6] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\m_blake2.m_hash256.m_matrix[9][17] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\m_blake2.m_hash256.m_matrix[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\m_blake2.m_hash256.v_q[0][31] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\m_blake2.m_hash256.v_q[0][7] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\m_blake2.m_hash256.v_q[3][4] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\m_blake2.m_hash256.v_q[0][22] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\m_io.m_config.ll_q[33] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\m_io.m_config.ll_q[45] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\m_blake2.m_hash256.m_matrix[12][21] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\m_blake2.m_hash256.m_matrix[12][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\m_blake2.m_hash256.v_q[0][1] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\m_io.m_config.ll_q[17] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\m_blake2.m_hash256.v_q[10][11] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\m_blake2.m_hash256.v_q[5][1] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\m_blake2.m_hash256.v_q[1][25] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\m_blake2.m_hash256.h_flat[19] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\m_blake2.m_hash256.m_matrix[9][25] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\m_blake2.m_hash256.v_q[4][28] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\m_io.m_config.ll_q[23] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\m_blake2.m_hash256.v_q[14][12] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\m_blake2.m_hash256.v_q[2][20] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\m_blake2.m_hash256.v_q[5][23] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\m_blake2.m_hash256.v_q[0][10] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\m_blake2.m_hash256.v_q[15][0] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\m_blake2.m_hash256.v_q[1][3] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\m_blake2.m_hash256.m_matrix[1][20] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\m_blake2.m_hash256.m_matrix[1][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\m_blake2.m_hash256.v_q[3][8] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[13] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\m_blake2.m_hash256.h_flat[29] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\m_blake2.m_hash256.v_q[14][30] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\m_blake2.m_hash256.v_q[2][29] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\m_blake2.m_hash256.v_q[5][3] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\m_blake2.m_hash256.h_flat[166] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\m_blake2.m_hash256.v_q[14][22] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\m_blake2.m_hash256.v_q[10][4] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\m_blake2.m_hash256.v_q[14][19] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\m_io.m_config.ll_q[0] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\m_blake2.m_hash256.v_q[13][28] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\m_blake2.m_hash256.v_q[1][8] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\m_blake2.m_hash256.v_q[4][0] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\m_blake2.m_hash256.v_q[14][14] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\m_blake2.m_hash256.v_q[6][7] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\m_blake2.m_hash256.v_q[6][25] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\m_blake2.m_hash256.m_matrix[1][26] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\m_blake2.m_hash256.v_q[1][29] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\m_blake2.m_hash256.v_q[6][17] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\m_blake2.m_hash256.m_matrix[3][31] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\m_blake2.m_hash256.v_q[6][2] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\m_blake2.m_hash256.v_q[6][13] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\m_blake2.m_hash256.v_q[2][2] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\m_blake2.m_hash256.v_q[6][12] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\m_blake2.m_hash256.v_q[0][15] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\m_blake2.m_hash256.v_q[5][29] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\m_blake2.m_hash256.m_matrix[8][21] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\m_blake2.m_hash256.m_matrix[8][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\m_blake2.m_hash256.round_q[5] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\m_blake2.m_hash256.round_q[6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\m_blake2.m_hash256.v_q[3][21] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\m_blake2.m_hash256.h_flat[150] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\m_blake2.m_hash256.v_q[0][30] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\m_blake2.m_hash256.m_matrix[5][31] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\m_blake2.m_hash256.m_matrix[5][5] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\m_blake2.m_hash256.v_q[4][4] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\m_blake2.m_hash256.v_q[0][21] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\m_blake2.m_hash256.v_q[9][21] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\m_blake2.m_hash256.v_q[5][9] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\m_blake2.m_hash256.v_q[6][16] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\m_blake2.m_hash256.m_matrix[11][6] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\m_blake2.m_hash256.m_matrix[10][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\m_blake2.m_hash256.v_q[0][19] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\m_blake2.m_hash256.m_matrix[12][25] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\m_blake2.m_hash256.m_matrix[12][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\m_blake2.m_hash256.v_q[5][21] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\m_blake2.m_hash256.v_q[6][8] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\m_blake2.m_hash256.v_q[1][1] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\m_blake2.m_hash256.v_q[10][16] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\m_blake2.m_hash256.v_q[11][20] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\m_blake2.m_hash256.v_q[3][25] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\m_blake2.m_hash256.v_q[5][17] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\m_blake2.m_hash256.h_flat[44] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\m_io.m_config.ll_q[34] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\m_blake2.m_hash256.m_matrix[1][12] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\m_blake2.m_hash256.v_q[2][4] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\m_blake2.m_hash256.h_flat[250] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\m_blake2.m_hash256.v_q[1][9] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\m_blake2.m_hash256.v_q[6][9] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\m_blake2.m_hash256.v_q[5][27] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\m_blake2.m_hash256.v_q[2][13] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\m_blake2.m_hash256.v_q[3][23] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\m_blake2.m_hash256.h_flat[124] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\m_blake2.m_hash256.v_q[4][1] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\m_blake2.m_hash256.m_matrix[12][18] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\m_blake2.m_hash256.v_q[5][18] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\m_blake2.m_hash256.v_q[11][24] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\m_blake2.m_hash256.v_q[10][29] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\m_blake2.m_hash256.v_q[3][20] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\m_blake2.m_hash256.v_q[0][25] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\m_blake2.m_hash256.h_flat[211] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\m_blake2.m_hash256.v_q[2][17] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\m_blake2.m_hash256.m_matrix[0][10] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\m_blake2.m_hash256.v_q[6][23] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\m_blake2.m_hash256.v_q[0][12] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\m_blake2.m_hash256.m_matrix[10][12] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\m_blake2.m_hash256.v_q[14][4] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\m_blake2.m_hash256.v_q[0][23] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\m_blake2.m_hash256.m_matrix[0][1] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\m_blake2.m_hash256.v_q[2][27] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\m_io.m_config.ll_q[15] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\m_blake2.m_hash256.v_q[2][5] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\m_blake2.m_hash256.v_q[9][25] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\m_blake2.m_hash256.v_q[1][10] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\m_blake2.m_hash256.v_q[1][4] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\m_blake2.m_hash256.v_q[2][23] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\m_blake2.m_hash256.v_q[5][13] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\m_blake2.m_hash256.v_q[3][27] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\m_blake2.m_hash256.h_flat[208] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\m_blake2.m_hash256.v_q[10][20] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\m_blake2.m_hash256.v_q[5][20] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\m_blake2.m_hash256.v_q[6][14] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\m_blake2.m_hash256.v_q[1][20] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\m_blake2.m_hash256.h_flat[194] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\m_blake2.m_hash256.v_q[6][24] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\m_blake2.m_hash256.v_q[0][14] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\m_blake2.m_hash256.v_q[11][28] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\m_blake2.m_hash256.v_q[5][15] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\m_blake2.m_hash256.v_q[2][30] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\m_blake2.m_hash256.v_q[1][23] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\m_blake2.m_hash256.v_q[2][9] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\m_blake2.m_hash256.v_q[9][12] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\m_blake2.m_hash256.m_matrix[0][26] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\m_blake2.m_hash256.m_matrix[0][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\m_blake2.m_hash256.v_q[15][24] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\m_blake2.m_hash256.m_matrix[0][12] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\m_io.m_config.ll_q[25] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\m_blake2.m_hash256.v_q[7][5] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\m_blake2.m_hash256.v_q[1][13] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\m_blake2.m_hash256.v_q[14][8] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\m_blake2.m_hash256.m_matrix[3][23] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\m_blake2.m_hash256.v_q[0][24] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\m_blake2.m_hash256.m_matrix[12][29] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\m_blake2.m_hash256.m_matrix[12][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\m_blake2.m_hash256.v_q[7][3] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\m_blake2.m_hash256.v_q[2][15] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\m_blake2.m_hash256.m_matrix[13][1] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\m_blake2.m_hash256.v_q[3][6] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\m_blake2.m_hash256.v_q[2][0] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\m_blake2.m_hash256.h_flat[198] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\m_blake2.m_hash256.v_q[1][14] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\m_blake2.m_hash256.v_q[0][0] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\m_blake2.m_hash256.m_matrix[11][11] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\m_blake2.m_hash256.v_q[3][28] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\m_io.m_config.ll_q[11] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\m_blake2.m_hash256.v_q[2][24] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\m_blake2.m_hash256.v_q[5][12] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\m_blake2.m_hash256.m_matrix[0][17] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\m_blake2.m_hash256.v_q[13][8] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\m_blake2.m_hash256.v_q[2][26] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\m_io.m_config.ll_q[60] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\m_blake2.m_hash256.v_q[15][18] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\m_blake2.m_hash256.m_matrix[6][21] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[16] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\m_blake2.m_hash256.m_matrix[14][28] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[24] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\m_blake2.m_hash256.v_q[5][19] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\m_blake2.m_hash256.v_q[3][0] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\m_blake2.m_hash256.v_q[14][26] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\m_blake2.m_hash256.m_matrix[7][19] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\m_blake2.m_hash256.m_matrix[7][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\m_blake2.m_hash256.m_matrix[11][26] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\m_blake2.m_hash256.m_matrix[11][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\m_blake2.m_hash256.v_q[2][1] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\m_blake2.m_hash256.v_q[6][11] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\m_blake2.m_hash256.v_q[12][11] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\m_blake2.m_hash256.v_q[3][29] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\m_io.m_config.ll_q[9] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\m_io.m_config.ll_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\m_blake2.m_hash256.m_matrix[14][26] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\m_blake2.m_hash256.m_matrix[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\m_blake2.m_hash256.v_q[15][28] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\m_blake2.m_hash256.v_q[2][19] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\m_blake2.m_hash256.v_q[15][12] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\m_blake2.m_hash256.v_q[15][6] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\m_blake2.m_hash256.m_matrix[4][27] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\m_blake2.m_hash256.m_matrix[4][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\m_blake2.m_hash256.v_q[14][31] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\m_blake2.m_hash256.m_matrix[8][3] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\m_blake2.m_hash256.m_matrix[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\m_blake2.m_hash256.m_matrix[10][15] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\m_blake2.m_hash256.m_matrix[10][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\m_blake2.m_hash256.m_matrix[2][12] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\m_blake2.m_hash256.m_matrix[2][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\m_blake2.m_hash256.v_q[5][24] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\m_blake2.m_hash256.v_q[4][5] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\m_blake2.m_hash256.v_q[13][14] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\m_blake2.m_hash256.v_q[5][22] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\m_blake2.m_hash256.m_matrix[15][20] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\m_blake2.m_hash256.v_q[5][30] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\m_blake2.m_hash256.m_matrix[6][13] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\m_blake2.m_hash256.m_matrix[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\m_blake2.m_hash256.m_matrix[1][17] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\m_blake2.m_hash256.m_matrix[1][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\m_blake2.m_hash256.v_q[7][6] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\m_blake2.m_hash256.v_q[1][16] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\m_blake2.m_hash256.v_q[1][19] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\m_blake2.m_hash256.m_matrix[8][31] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\m_blake2.m_hash256.m_matrix[8][31]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\m_blake2.m_hash256.v_q[15][27] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\m_blake2.m_hash256.v_q[1][5] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\m_blake2.m_hash256.v_q[2][31] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\m_blake2.m_hash256.m_matrix[3][2] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\m_blake2.m_hash256.m_matrix[8][22] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\m_blake2.m_hash256.m_matrix[8][14]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\m_blake2.m_hash256.m_matrix[7][15] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\m_blake2.m_hash256.v_q[7][18] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\m_blake2.m_hash256.v_q[6][15] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\m_blake2.m_hash256.v_q[6][29] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\m_blake2.m_hash256.v_q[2][6] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\m_blake2.m_hash256.m_matrix[2][26] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\m_blake2.m_hash256.v_q[15][16] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\m_io.m_config.ll_q[26] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\m_blake2.m_hash256.m_matrix[14][5] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\m_blake2.m_hash256.v_q[8][30] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\m_blake2.m_hash256.v_q[10][12] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\m_blake2.m_hash256.m_matrix[8][26] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\m_blake2.m_hash256.v_q[15][25] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\m_blake2.m_hash256.v_q[9][5] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\m_blake2.m_hash256.v_q[5][10] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\m_blake2.m_hash256.m_matrix[11][3] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\m_blake2.m_hash256.m_matrix[5][8] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\m_blake2.m_hash256.v_q[15][2] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\m_blake2.m_hash256.v_q[6][20] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\m_blake2.m_hash256.m_matrix[9][23] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\m_blake2.m_hash256.m_matrix[9][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\m_blake2.m_hash256.v_q[7][22] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\m_blake2.m_hash256.v_q[2][25] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\m_blake2.m_hash256.m_matrix[9][3] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\m_blake2.m_hash256.m_matrix[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\m_blake2.m_hash256.v_q[1][24] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\m_blake2.m_hash256.v_q[5][0] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\m_blake2.m_hash256.v_q[7][11] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\m_blake2.m_hash256.v_q[7][1] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\m_blake2.m_hash256.v_q[15][26] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\m_blake2.m_hash256.v_q[3][22] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\m_blake2.m_hash256.v_q[8][21] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\m_blake2.m_hash256.v_q[10][30] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\m_blake2.m_hash256.v_q[1][31] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\m_blake2.m_hash256.h_flat[28] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\m_blake2.m_hash256.m_matrix[7][0] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\m_blake2.m_hash256.m_matrix[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\m_blake2.m_hash256.v_q[14][11] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\m_blake2.m_hash256.v_q[5][14] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\m_io.m_config.ll_q[50] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\m_blake2.m_hash256.m_matrix[7][26] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\m_blake2.m_hash256.m_matrix[7][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\m_blake2.m_hash256.v_q[3][3] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\m_blake2.m_hash256.m_matrix[12][27] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\m_blake2.m_hash256.v_q[7][27] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\m_blake2.m_hash256.v_q[3][26] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\m_blake2.m_hash256.v_q[13][22] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\m_blake2.m_hash256.m_matrix[11][14] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\m_io.m_config.ll_q[51] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\m_blake2.m_hash256.h_flat[179] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\m_blake2.m_hash256.v_q[3][15] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\m_blake2.m_hash256.v_q[11][8] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\m_blake2.m_hash256.v_q[1][21] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\m_blake2.m_hash256.v_q[0][8] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\m_blake2.m_hash256.m_matrix[4][23] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\m_blake2.m_hash256.m_matrix[11][1] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\m_blake2.m_hash256.m_matrix[10][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\m_blake2.m_hash256.v_q[5][6] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\m_blake2.m_hash256.m_matrix[4][18] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\m_blake2.m_hash256.m_matrix[4][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\m_blake2.m_hash256.m_matrix[2][4] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\m_blake2.m_hash256.v_q[7][30] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\m_blake2.m_hash256.v_q[10][2] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\m_blake2.m_hash256.m_matrix[10][28] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\m_blake2.m_hash256.m_matrix[10][11] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\m_blake2.m_hash256.m_matrix[10][27] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\m_blake2.m_hash256.h_flat[144] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\m_blake2.m_hash256.v_q[1][18] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\m_blake2.m_hash256.m_matrix[8][7] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\m_blake2.m_hash256.m_matrix[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\m_blake2.m_hash256.v_q[12][18] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\m_blake2.m_hash256.v_q[0][29] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\m_blake2.m_hash256.m_matrix[5][26] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\m_blake2.m_hash256.m_matrix[5][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\m_blake2.m_hash256.v_q[11][29] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\m_blake2.m_hash256.m_matrix[2][18] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\m_io.m_config.ll_q[48] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\m_io.m_config.ll_q[31] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\m_blake2.m_hash256.v_q[1][26] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\m_blake2.m_hash256.v_q[7][0] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\m_blake2.m_hash256.m_matrix[8][17] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\m_blake2.m_hash256.m_matrix[8][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\m_blake2.m_hash256.m_matrix[15][21] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\m_blake2.m_hash256.m_matrix[11][10] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\m_blake2.m_hash256.m_matrix[11][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\m_blake2.m_hash256.h_flat[159] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\m_io.m_config.cfg_cnt_q[3] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\m_blake2.m_hash256.v_q[3][7] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\m_blake2.m_hash256.m_matrix[11][22] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\m_blake2.m_hash256.v_q[0][2] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\m_blake2.m_hash256.m_matrix[10][10] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\m_blake2.m_hash256.m_matrix[10][10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\m_blake2.m_hash256.m_matrix[13][17] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\m_blake2.m_hash256.m_matrix[13][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\m_blake2.m_hash256.v_q[15][1] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\m_blake2.m_hash256.v_q[7][7] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\m_blake2.m_hash256.m_matrix[7][31] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\m_blake2.m_hash256.v_q[2][12] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\m_blake2.m_hash256.v_q[14][24] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\m_blake2.m_hash256.v_q[10][24] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\m_blake2.m_hash256.v_q[2][21] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\m_blake2.m_hash256.m_matrix[10][7] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\m_blake2.m_hash256.m_matrix[4][26] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\m_blake2.m_hash256.m_matrix[4][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\m_blake2.m_hash256.v_q[7][4] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\m_blake2.m_hash256.v_q[10][6] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\m_blake2.m_hash256.v_q[14][0] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\m_blake2.m_hash256.v_q[5][7] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\m_blake2.m_hash256.v_q[9][29] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\m_blake2.m_hash256.m_matrix[0][22] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\m_blake2.m_hash256.v_q[2][3] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\m_blake2.m_hash256.v_q[1][6] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\m_blake2.m_hash256.v_q[1][22] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\m_blake2.m_hash256.v_q[15][11] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\m_blake2.m_hash256.m_matrix[9][15] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\m_blake2.m_hash256.v_q[3][14] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\m_blake2.m_hash256.v_q[8][13] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\m_blake2.m_hash256.m_matrix[0][11] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\m_blake2.m_hash256.m_matrix[0][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\m_blake2.m_hash256.v_q[15][14] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\m_blake2.m_hash256.v_q[12][26] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\m_blake2.m_hash256.v_q[15][15] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\m_blake2.m_hash256.v_q[3][13] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\m_blake2.m_hash256.v_q[10][25] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\m_blake2.m_hash256.m_matrix[5][24] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\m_blake2.m_hash256.m_matrix[5][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\m_blake2.m_hash256.v_q[3][19] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\m_blake2.m_hash256.m_matrix[1][9] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\m_blake2.m_hash256.v_q[9][8] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\m_blake2.m_hash256.v_q[11][11] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\m_blake2.m_hash256.m_matrix[9][1] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\m_blake2.m_hash256.m_matrix[8][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\m_blake2.m_hash256.m_matrix[3][26] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\m_blake2.m_hash256.m_matrix[3][26]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\m_blake2.m_hash256.m_matrix[5][20] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\m_blake2.m_hash256.m_matrix[5][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\m_blake2.m_hash256.m_matrix[8][30] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\m_blake2.m_hash256.v_q[4][24] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\m_blake2.m_hash256.v_q[3][1] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\m_blake2.m_hash256.m_matrix[2][10] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\m_blake2.m_hash256.m_matrix[11][9] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\m_blake2.m_hash256.v_q[1][28] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\m_blake2.m_hash256.m_matrix[12][26] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\m_blake2.m_hash256.v_q[3][31] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\m_blake2.m_hash256.v_q[8][10] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\m_blake2.m_hash256.v_q[1][27] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\m_blake2.m_hash256.v_q[7][31] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\m_blake2.m_hash256.h_flat[253] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\m_blake2.m_hash256.v_q[12][19] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\m_blake2.m_hash256.v_q[1][15] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\m_blake2.m_hash256.v_q[10][5] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\m_blake2.m_hash256.v_q[14][6] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\m_blake2.m_hash256.m_matrix[2][3] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\m_blake2.m_hash256.m_matrix[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\m_blake2.m_hash256.m_matrix[15][12] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\m_blake2.m_hash256.v_q[9][16] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\m_blake2.m_hash256.m_matrix[6][19] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\m_blake2.m_hash256.m_matrix[6][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\m_blake2.m_hash256.v_q[13][2] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\m_blake2.m_hash256.m_matrix[2][2] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\m_blake2.m_hash256.v_q[8][11] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\m_blake2.m_hash256.m_matrix[2][23] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\m_blake2.m_hash256.m_matrix[2][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\m_blake2.m_hash256.m_matrix[3][27] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\m_blake2.m_hash256.v_q[8][8] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\m_blake2.m_hash256.v_q[14][10] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\m_blake2.m_hash256.m_matrix[11][17] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\m_blake2.m_hash256.m_matrix[11][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\m_blake2.m_hash256.v_q[2][10] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\m_blake2.m_hash256.v_q[2][8] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\m_blake2.m_hash256.m_matrix[5][23] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\m_blake2.m_hash256.v_q[13][18] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\m_blake2.m_hash256.v_q[12][27] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\m_blake2.m_hash256.m_matrix[8][9] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\m_blake2.m_hash256.v_q[3][16] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\m_blake2.m_hash256.h_flat[243] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\m_blake2.m_hash256.v_q[10][13] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\m_blake2.m_hash256.v_q[9][0] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\m_blake2.m_hash256.m_matrix[10][22] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\m_blake2.m_hash256.m_matrix[10][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\m_blake2.m_hash256.h_flat[220] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\m_blake2.m_hash256.m_matrix[9][7] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\m_blake2.m_hash256.m_matrix[13][6] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\m_blake2.m_hash256.m_matrix[5][18] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\m_blake2.m_hash256.m_matrix[9][31] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\m_blake2.m_hash256.v_q[3][30] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\m_blake2.m_hash256.m_matrix[15][17] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\m_blake2.m_hash256.v_q[15][23] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\m_blake2.m_hash256.v_q[3][2] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\m_blake2.m_hash256.v_q[7][21] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\m_blake2.m_hash256.v_q[5][16] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\m_blake2.m_hash256.m_matrix[1][27] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\m_blake2.m_hash256.m_matrix[7][11] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\m_blake2.m_hash256.v_q[8][25] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\m_blake2.m_hash256.v_q[11][12] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\m_blake2.m_hash256.v_q[2][28] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\m_blake2.m_hash256.m_matrix[3][28] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\m_blake2.m_hash256.v_q[8][6] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\m_blake2.m_hash256.m_matrix[10][1] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\m_blake2.m_hash256.m_matrix[10][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\m_blake2.m_hash256.m_matrix[3][18] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\m_blake2.m_hash256.v_q[2][22] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\m_blake2.m_hash256.m_matrix[5][12] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\m_blake2.m_hash256.v_q[1][12] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\m_blake2.m_hash256.v_q[0][4] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\m_blake2.m_hash256.m_matrix[14][20] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\m_blake2.m_hash256.m_matrix[1][11] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\m_blake2.m_hash256.m_matrix[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\m_blake2.m_hash256.v_q[6][19] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\m_blake2.m_hash256.v_q[8][3] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\m_blake2.m_hash256.v_q[10][8] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\m_blake2.m_hash256.v_q[13][0] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\m_blake2.m_hash256.m_matrix[5][28] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\m_blake2.m_hash256.v_q[0][9] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\m_blake2.m_hash256.m_matrix[7][14] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\m_blake2.m_hash256.m_matrix[6][0] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\m_blake2.m_hash256.m_matrix[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\m_blake2.m_hash256.m_matrix[6][12] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\m_blake2.m_hash256.m_matrix[9][22] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\m_blake2.m_hash256.m_matrix[9][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\m_blake2.m_hash256.m_matrix[13][9] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\m_blake2.m_hash256.v_q[8][15] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\m_blake2.m_hash256.v_q[7][23] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\m_blake2.m_hash256.v_q[1][7] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\m_blake2.m_hash256.m_matrix[8][27] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\m_blake2.m_hash256.v_q[3][5] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\m_blake2.m_hash256.v_q[1][30] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\m_blake2.m_hash256.v_q[8][12] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\m_blake2.m_hash256.m_matrix[5][16] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\m_blake2.m_hash256.v_q[11][3] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\m_blake2.m_hash256.v_q[7][9] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\m_io.m_config.ll_q[35] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\m_blake2.m_hash256.m_matrix[5][0] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\m_blake2.m_hash256.v_q[5][26] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\m_blake2.m_hash256.v_q[15][20] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\m_blake2.m_hash256.v_q[7][26] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\m_blake2.m_hash256.m_matrix[0][19] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\m_blake2.m_hash256.m_matrix[13][29] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\m_blake2.m_hash256.v_q[7][19] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\m_blake2.m_hash256.v_q[7][8] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\m_blake2.m_hash256.v_q[15][19] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\m_blake2.m_hash256.v_q[15][31] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\m_blake2.m_hash256.v_q[13][10] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\m_blake2.m_hash256.v_q[13][3] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\m_blake2.m_hash256.h_flat[32] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\m_blake2.m_hash256.m_matrix[2][19] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\m_blake2.m_hash256.m_matrix[2][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\m_blake2.m_hash256.v_q[15][4] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\m_blake2.m_hash256.m_matrix[15][19] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\m_blake2.m_hash256.m_matrix[15][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\m_blake2.m_hash256.v_q[15][3] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\m_blake2.m_hash256.m_matrix[9][20] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\m_blake2.m_hash256.m_matrix[9][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\m_blake2.m_hash256.v_q[8][22] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\m_blake2.m_hash256.m_matrix[7][2] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\m_blake2.m_hash256.m_matrix[7][27] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\m_blake2.m_hash256.v_q[14][2] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\m_blake2.m_hash256.v_q[14][28] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\m_blake2.m_hash256.v_q[7][12] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\m_blake2.m_hash256.v_q[11][13] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\m_blake2.m_hash256.m_matrix[1][15] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\m_blake2.m_hash256.v_q[8][20] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\m_blake2.m_hash256.v_q[6][28] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[4] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[56] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\m_blake2.m_hash256.v_q[12][5] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\m_blake2.m_hash256.v_q[0][13] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\m_blake2.m_hash256.h_flat[214] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\m_blake2.m_hash256.v_q[8][29] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\m_blake2.m_hash256.v_q[8][24] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\m_blake2.m_hash256.v_q[7][13] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\m_blake2.m_hash256.v_q[8][18] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\m_blake2.m_hash256.v_q[3][12] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\m_blake2.m_hash256.m_matrix[4][10] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\m_blake2.m_hash256.m_matrix[15][13] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\m_blake2.m_hash256.m_matrix[9][11] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\m_blake2.m_hash256.m_matrix[9][11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\m_blake2.m_hash256.v_q[2][7] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\m_blake2.m_hash256.v_q[8][5] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\m_blake2.m_hash256.m_matrix[11][20] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\m_blake2.m_hash256.m_matrix[11][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\m_blake2.m_hash256.m_matrix[8][24] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\m_blake2.m_hash256.m_matrix[8][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\m_blake2.m_hash256.m_matrix[2][17] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\m_blake2.m_hash256.m_matrix[2][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\m_blake2.m_hash256.v_q[12][10] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\m_blake2.m_hash256.m_matrix[0][14] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\m_blake2.m_hash256.m_matrix[5][6] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\m_blake2.m_hash256.m_matrix[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\m_blake2.m_hash256.v_q[7][20] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\m_blake2.m_hash256.m_matrix[8][13] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\m_blake2.m_hash256.m_matrix[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\m_blake2.m_hash256.v_q[12][24] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\m_blake2.m_hash256.v_q[9][11] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\m_blake2.m_hash256.v_q[7][17] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\m_blake2.m_hash256.m_matrix[13][24] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\m_blake2.m_hash256.v_q[7][2] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\m_blake2.m_hash256.m_matrix[4][2] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\m_blake2.m_hash256.h_flat[25] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\m_blake2.m_hash256.m_matrix[1][8] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\m_blake2.m_hash256.m_matrix[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\m_blake2.m_hash256.m_matrix[15][6] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\m_blake2.m_hash256.m_matrix[15][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\m_blake2.m_hash256.v_q[13][30] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\m_blake2.m_hash256.v_q[7][10] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\m_blake2.m_hash256.m_matrix[13][21] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\m_blake2.m_hash256.v_q[11][4] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\m_blake2.m_hash256.m_matrix[2][11] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\m_blake2.m_hash256.v_q[15][21] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\m_blake2.m_hash256.v_q[7][16] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\m_blake2.m_hash256.m_matrix[13][16] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\m_blake2.m_hash256.m_matrix[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\m_blake2.m_hash256.v_q[0][11] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\m_blake2.m_hash256.v_q[8][7] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\m_blake2.m_hash256.m_matrix[9][12] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\m_blake2.m_hash256.m_matrix[3][0] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\m_blake2.m_hash256.m_matrix[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\m_blake2.m_hash256.m_matrix[4][5] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\m_blake2.m_hash256.m_matrix[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\m_blake2.m_hash256.m_matrix[1][13] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\m_blake2.m_hash256.m_matrix[15][23] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\m_blake2.m_hash256.v_q[9][13] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\m_blake2.m_hash256.v_q[7][14] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\m_blake2.m_hash256.m_matrix[8][6] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\m_blake2.m_hash256.m_matrix[5][4] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\m_blake2.m_hash256.m_matrix[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\m_blake2.m_hash256.v_q[10][22] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\m_blake2.m_hash256.m_matrix[1][4] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\m_blake2.m_hash256.m_matrix[0][21] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\m_blake2.m_hash256.m_matrix[0][21]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\m_blake2.m_hash256.m_matrix[10][14] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\m_blake2.m_hash256.m_matrix[1][7] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\m_blake2.m_hash256.m_matrix[5][19] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\m_blake2.m_hash256.m_matrix[5][19]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\m_blake2.m_hash256.m_matrix[4][28] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\m_blake2.m_hash256.v_q[8][19] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\m_blake2.m_hash256.m_matrix[1][16] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\m_blake2.m_hash256.m_matrix[1][16]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\m_blake2.m_hash256.v_q[9][14] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\m_blake2.m_hash256.v_q[9][4] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\m_blake2.m_hash256.v_q[12][28] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\m_blake2.m_hash256.v_q[12][0] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\m_blake2.m_hash256.v_q[11][10] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\m_blake2.m_hash256.m_matrix[0][15] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\m_blake2.m_hash256.m_matrix[0][15]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\m_blake2.m_hash256.m_matrix[6][26] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\m_blake2.m_hash256.m_matrix[10][17] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\m_blake2.m_hash256.m_matrix[10][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\m_blake2.m_hash256.m_matrix[2][8] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\m_blake2.m_hash256.v_q[13][16] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\m_blake2.m_hash256.v_q[11][17] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\m_blake2.m_hash256.m_matrix[2][15] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\m_blake2.m_hash256.m_matrix[5][29] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\m_blake2.m_hash256.m_matrix[5][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\m_blake2.m_hash256.m_matrix[2][13] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\m_blake2.m_hash256.h_flat[230] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\m_blake2.m_hash256.v_q[7][29] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\m_blake2.m_hash256.m_matrix[7][30] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\m_blake2.m_hash256.m_matrix[3][24] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\m_blake2.m_hash256.m_matrix[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\m_blake2.m_hash256.m_matrix[12][0] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\m_blake2.m_hash256.v_q[11][1] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\m_blake2.m_hash256.h_flat[172] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\m_blake2.m_hash256.m_matrix[6][18] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\m_blake2.m_hash256.m_matrix[6][2] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\m_blake2.m_hash256.m_matrix[5][10] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\m_blake2.m_hash256.v_q[13][6] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\m_blake2.m_hash256.m_matrix[4][29] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\m_blake2.m_hash256.m_matrix[7][4] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\m_blake2.m_hash256.m_matrix[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\m_blake2.m_hash256.m_matrix[2][24] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\m_blake2.m_hash256.m_matrix[3][12] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\m_blake2.m_hash256.m_matrix[9][19] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\m_blake2.m_hash256.m_matrix[14][31] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\m_blake2.m_hash256.v_q[14][25] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\m_blake2.m_hash256.v_q[8][26] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\m_blake2.m_hash256.v_q[13][26] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\m_blake2.m_hash256.m_matrix[4][30] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\m_blake2.m_hash256.m_matrix[7][8] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\m_blake2.m_hash256.m_matrix[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\m_blake2.m_hash256.m_matrix[4][21] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\m_blake2.m_hash256.m_matrix[1][19] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\m_blake2.m_hash256.m_matrix[15][2] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\m_blake2.m_hash256.v_q[11][0] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\m_blake2.m_hash256.m_matrix[8][15] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\m_blake2.m_hash256.v_q[8][28] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\m_blake2.m_hash256.m_matrix[12][17] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\m_blake2.m_hash256.m_matrix[12][9]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\m_blake2.m_hash256.m_matrix[3][19] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\m_blake2.m_hash256.m_matrix[12][8] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\m_blake2.m_hash256.v_q[6][31] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\m_blake2.m_hash256.m_matrix[3][29] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\m_blake2.m_hash256.m_matrix[4][24] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\m_blake2.m_hash256.m_matrix[13][13] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\m_blake2.m_hash256.h_flat[112] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\m_blake2.m_hash256.v_q[14][3] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\m_blake2.m_hash256.m_matrix[10][21] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\m_blake2.m_hash256.v_q[12][12] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\m_blake2.m_hash256.v_q[7][28] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\m_blake2.m_hash256.v_q[12][20] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\m_blake2.m_hash256.v_q[8][0] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\m_blake2.m_hash256.m_matrix[4][16] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\m_blake2.m_hash256.m_matrix[1][28] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\m_blake2.m_hash256.m_matrix[2][22] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\m_blake2.m_hash256.m_matrix[2][27] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\m_blake2.m_hash256.v_q[8][4] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\m_blake2.m_hash256.v_q[7][25] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\m_blake2.m_hash256.v_q[14][18] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\m_blake2.m_hash256.m_matrix[5][2] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\m_blake2.m_hash256.m_matrix[3][21] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\m_blake2.m_hash256.m_matrix[1][2] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\m_blake2.m_hash256.m_matrix[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\m_blake2.m_hash256.v_q[13][20] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\m_blake2.m_hash256.v_q[11][22] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\m_blake2.m_hash256.m_matrix[7][12] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\m_blake2.m_hash256.m_matrix[7][12]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\m_blake2.m_hash256.v_q[5][8] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\m_blake2.m_hash256.m_matrix[8][19] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\m_blake2.m_hash256.m_matrix[4][6] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\m_blake2.m_hash256.m_matrix[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\m_io.m_config.ll_q[24] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\m_blake2.m_hash256.v_q[13][19] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\m_blake2.m_hash256.m_matrix[4][8] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\m_blake2.m_hash256.m_matrix[11][29] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\m_blake2.m_hash256.m_matrix[11][29]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\m_blake2.m_hash256.v_q[11][30] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\m_blake2.m_hash256.m_matrix[6][27] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\m_blake2.m_hash256.m_matrix[6][27]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\m_blake2.m_hash256.m_matrix[10][9] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\m_blake2.m_hash256.m_matrix[8][11] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\m_blake2.m_hash256.v_q[10][15] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\m_blake2.m_hash256.v_q[12][2] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\m_blake2.m_hash256.m_matrix[7][17] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\m_blake2.m_hash256.v_q[9][6] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\m_blake2.m_hash256.m_matrix[3][22] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\m_blake2.m_hash256.m_matrix[1][0] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\m_blake2.m_hash256.m_matrix[3][30] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\m_blake2.m_hash256.m_matrix[3][4] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\m_blake2.m_hash256.m_matrix[0][16] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\m_blake2.m_hash256.m_matrix[3][11] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\m_blake2.m_hash256.m_matrix[15][15] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\m_blake2.m_hash256.m_matrix[7][3] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[40] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\m_blake2.m_hash256.m_matrix[2][30] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\m_blake2.m_hash256.m_matrix[2][22]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\m_blake2.m_hash256.m_matrix[13][5] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\m_blake2.m_hash256.h_flat[64] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\m_blake2.m_hash256.v_q[9][22] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\m_blake2.m_hash256.v_q[2][18] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\m_blake2.m_hash256.m_matrix[3][15] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\m_blake2.m_hash256.m_matrix[4][22] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\m_blake2.m_hash256.v_q[4][12] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\m_blake2.m_hash256.v_q[12][9] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\m_blake2.m_hash256.v_q[15][17] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\m_blake2.m_hash256.m_matrix[5][22] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\m_blake2.m_hash256.v_q[11][14] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\m_blake2.m_hash256.h_flat[246] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\m_blake2.m_hash256.v_q[13][11] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\m_blake2.m_hash256.v_q[13][27] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\m_blake2.m_hash256.m_matrix[10][13] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\m_blake2.m_hash256.m_matrix[3][13] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\m_blake2.m_hash256.m_matrix[7][20] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\m_blake2.m_hash256.m_matrix[7][20]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\m_blake2.m_hash256.m_matrix[13][19] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\m_blake2.m_hash256.v_q[10][19] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\m_blake2.m_hash256.m_matrix[12][16] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\m_blake2.m_hash256.m_matrix[3][16] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\m_blake2.m_hash256.m_matrix[6][25] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\m_blake2.m_hash256.v_q[15][7] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\m_blake2.m_hash256.v_q[8][14] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\m_blake2.m_hash256.m_matrix[13][27] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\m_blake2.m_hash256.v_q[9][30] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\m_blake2.m_hash256.m_matrix[3][7] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\m_blake2.m_hash256.m_matrix[12][11] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\m_blake2.m_hash256.m_matrix[11][5] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\m_blake2.m_hash256.m_matrix[1][6] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\m_io.m_config.ll_q[43] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\m_blake2.m_hash256.v_q[14][17] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\m_blake2.m_hash256.v_q[9][17] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\m_blake2.m_hash256.m_matrix[7][21] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\m_blake2.m_hash256.v_q[11][21] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\data[5] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\m_blake2.m_hash256.v_q[12][3] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\m_blake2.m_hash256.m_matrix[9][6] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\m_blake2.m_hash256.m_matrix[3][5] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\m_blake2.m_hash256.m_matrix[6][28] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[22] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\m_blake2.m_hash256.m_matrix[13][22] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\m_blake2.m_hash256.res_cnt_q[5] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\m_blake2.m_hash256.v_q[15][5] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\m_blake2.m_hash256.m_matrix[7][16] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\m_blake2.m_hash256.m_matrix[3][17] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\m_blake2.m_hash256.m_matrix[14][8] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\m_blake2.m_hash256.m_matrix[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\m_blake2.m_hash256.m_matrix[3][3] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\m_blake2.m_hash256.h_flat[160] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\m_blake2.m_hash256.v_q[11][26] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\m_blake2.m_hash256.m_matrix[11][7] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\m_io.m_config.ll_q[28] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\m_blake2.m_hash256.m_matrix[14][21] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\m_blake2.m_hash256.m_matrix[2][29] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\m_blake2.m_hash256.m_matrix[8][16] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\m_blake2.m_hash256.m_matrix[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\m_blake2.m_hash256.v_q[7][24] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\m_blake2.m_hash256.m_matrix[5][14] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\m_blake2.m_hash256.m_matrix[14][6] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\m_blake2.m_hash256.m_matrix[14][24] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\m_blake2.m_hash256.m_matrix[7][22] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\m_blake2.m_hash256.m_matrix[14][1] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\m_blake2.m_hash256.fsm_q[2] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\m_blake2.m_hash256.m_matrix[10][18] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\m_blake2.m_hash256.v_q[10][0] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\m_blake2.m_hash256.m_matrix[4][13] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\m_blake2.m_hash256.m_matrix[4][20] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\m_blake2.m_hash256.m_matrix[5][7] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\m_blake2.m_hash256.m_matrix[4][14] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\m_blake2.m_hash256.m_matrix[14][2] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\m_blake2.m_hash256.v_q[12][16] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\m_blake2.m_hash256.m_matrix[6][14] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\m_blake2.m_hash256.m_matrix[5][30] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\m_blake2.m_hash256.v_q[9][7] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\m_blake2.m_hash256.v_q[9][10] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\m_blake2.m_hash256.m_matrix[1][24] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\m_blake2.m_hash256.v_q[9][3] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\m_blake2.m_hash256.m_matrix[12][3] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\m_blake2.m_hash256.v_q[8][31] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\m_blake2.m_hash256.v_q[14][7] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\m_blake2.m_hash256.m_matrix[6][11] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\m_blake2.m_hash256.m_matrix[4][17] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\m_blake2.m_hash256.m_matrix[2][9] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\m_blake2.m_hash256.m_matrix[2][25] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\m_blake2.m_hash256.m_matrix[14][18] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(\m_blake2.m_hash256.v_q[15][13] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\m_blake2.m_hash256.m_matrix[13][26] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\m_blake2.m_hash256.v_q[11][25] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\m_blake2.m_hash256.m_matrix[2][5] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\m_blake2.m_hash256.h_flat[88] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\m_blake2.m_hash256.m_matrix[12][9] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\m_blake2.m_hash256.m_matrix[12][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\m_io.m_config.ll_q[19] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\m_io.m_config.ll_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\m_blake2.m_hash256.v_q[11][5] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\m_blake2.m_hash256.m_matrix[4][12] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\m_io.m_config.kk_q[1] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\m_blake2.m_hash256.v_q[10][17] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\m_blake2.m_hash256.m_matrix[6][3] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\m_blake2.m_hash256.m_matrix[14][22] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\m_blake2.m_hash256.m_matrix[11][21] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\m_blake2.m_hash256.v_q[14][29] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\m_blake2.m_hash256.m_matrix[4][25] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\m_blake2.m_hash256.m_matrix[4][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\m_blake2.m_hash256.m_matrix[13][25] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\m_blake2.m_hash256.v_q[9][1] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\m_blake2.m_hash256.m_matrix[9][30] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\m_blake2.m_hash256.m_matrix[6][9] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\m_blake2.m_hash256.m_matrix[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\m_blake2.m_hash256.m_matrix[12][20] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\m_blake2.m_hash256.m_matrix[8][28] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\m_blake2.m_hash256.m_matrix[8][28]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\m_blake2.m_hash256.m_matrix[11][31] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\m_blake2.m_hash256.m_matrix[11][23]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\m_blake2.m_hash256.v_q[11][6] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\m_blake2.m_hash256.v_q[12][8] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\m_blake2.m_hash256.v_q[9][19] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\m_blake2.m_hash256.m_matrix[14][16] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\m_blake2.m_hash256.m_matrix[8][0] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\m_blake2.m_hash256.m_matrix[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\m_blake2.m_hash256.m_matrix[2][1] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(\m_blake2.m_hash256.m_matrix[2][20] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\m_blake2.m_hash256.v_q[12][6] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\m_blake2.m_hash256.m_matrix[8][20] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\m_blake2.m_hash256.v_q[10][23] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\m_blake2.m_hash256.v_q[9][2] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\m_blake2.m_hash256.v_q[2][16] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\m_blake2.m_hash256.m_matrix[9][8] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\m_blake2.m_hash256.m_matrix[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(\m_blake2.m_hash256.v_q[10][10] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\m_io.m_config.ll_q[18] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\m_io.m_config.ll_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\m_blake2.m_hash256.v_q[12][22] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\m_blake2.m_hash256.m_matrix[7][5] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\m_blake2.m_hash256.m_matrix[9][16] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\m_blake2.m_hash256.v_q[12][14] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\m_blake2.m_hash256.m_matrix[3][8] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\m_blake2.m_hash256.v_q[14][9] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\m_blake2.m_hash256.m_matrix[4][1] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\m_blake2.m_hash256.m_matrix[12][28] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\m_blake2.m_hash256.m_matrix[3][1] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\m_blake2.m_hash256.m_matrix[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\m_blake2.m_hash256.m_matrix[13][7] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\m_blake2.m_hash256.m_matrix[12][5] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\m_blake2.m_hash256.v_q[7][15] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\m_blake2.m_hash256.m_matrix[13][18] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\m_blake2.m_hash256.m_matrix[13][18]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[46] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[44] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\m_blake2.m_hash256.m_matrix[0][29] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\m_blake2.m_hash256.v_q[12][25] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\m_blake2.m_hash256.m_matrix[15][1] ),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\m_blake2.m_hash256.m_matrix[9][4] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\m_blake2.m_hash256.v_q[11][16] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\m_blake2.m_hash256.m_matrix[10][0] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(\m_blake2.m_hash256.m_matrix[10][0]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\m_blake2.m_hash256.m_matrix[13][11] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(\m_blake2.m_hash256.m_matrix[12][1] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\m_blake2.m_hash256.m_matrix[11][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(\m_blake2.m_hash256.m_matrix[9][13] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\m_blake2.m_hash256.m_matrix[9][13]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(\m_blake2.m_hash256.v_q[15][29] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\m_blake2.m_hash256.m_matrix[11][28] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\m_blake2.m_hash256.m_matrix[12][22] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\m_blake2.m_hash256.m_matrix[5][3] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\m_blake2.m_hash256.m_matrix[2][31] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\m_blake2.m_hash256.m_matrix[8][2] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\m_blake2.m_hash256.round_q[0] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\m_blake2.m_hash256.v_q[13][25] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(\m_blake2.m_hash256.v_q[11][31] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\m_blake2.m_hash256.m_matrix[5][17] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(\m_blake2.m_hash256.m_matrix[5][17]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\m_blake2.m_hash256.v_q[10][3] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(\m_blake2.m_hash256.m_matrix[14][27] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\m_blake2.m_hash256.m_matrix[10][8] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(\m_blake2.m_hash256.m_matrix[9][21] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\m_blake2.m_hash256.h_flat[188] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(\m_blake2.m_hash256.v_q[15][9] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\m_blake2.m_hash256.v_q[8][27] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(\m_blake2.m_hash256.m_matrix[1][25] ),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\m_blake2.m_hash256.m_matrix[4][0] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(\m_blake2.m_hash256.v_q[12][1] ),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\m_blake2.m_hash256.m_matrix[5][27] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\m_blake2.m_hash256.m_matrix[9][28] ),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\m_blake2.m_hash256.m_matrix[13][10] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(\m_blake2.m_hash256.m_matrix[3][9] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\m_blake2.m_hash256.m_matrix[13][31] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(\m_blake2.m_hash256.m_matrix[7][1] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\m_blake2.m_hash256.m_matrix[15][14] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(\m_blake2.m_hash256.m_matrix[1][29] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\m_blake2.m_hash256.v_q[8][16] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(\m_blake2.m_hash256.m_matrix[3][6] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\m_blake2.m_hash256.m_matrix[2][30]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\m_blake2.m_hash256.m_matrix[12][6] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\m_blake2.m_hash256.v_q[13][17] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\m_blake2.m_hash256.m_matrix[7][28] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\m_blake2.m_hash256.m_matrix[6][16] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\m_blake2.m_hash256.v_q[12][30] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\m_blake2.m_hash256.m_matrix[5][9] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\m_blake2.m_hash256.v_q[4][3] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\m_blake2.m_hash256.m_matrix[9][18] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\m_blake2.m_hash256.v_q[11][2] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\m_blake2.m_hash256.m_matrix[9][10] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\m_blake2.m_hash256.v_q[8][1] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\m_io.m_config.cfg_cnt_q[2] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\m_blake2.m_hash256.v_q[13][9] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\m_blake2.m_hash256.v_q[13][31] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\m_blake2.m_hash256.v_q[8][2] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\m_blake2.m_hash256.h_flat[252] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\m_blake2.m_hash256.m_matrix[5][1] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\m_blake2.m_hash256.m_matrix[11][23] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[3] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\m_blake2.m_hash256.v_q[13][4] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(\m_blake2.m_hash256.v_q[12][17] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\m_blake2.m_hash256.m_matrix[12][31] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\m_blake2.m_hash256.v_q[9][31] ),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\m_blake2.m_hash256.m_matrix[2][28] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\m_blake2.m_hash256.v_q[8][23] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\m_blake2.m_hash256.m_matrix[12][4] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(\m_blake2.m_hash256.v_q[11][19] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\m_blake2.m_hash256.m_matrix[0][23] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(\m_blake2.m_hash256.v_q[12][29] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\m_io.m_config.ll_q[36] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(\m_blake2.m_hash256.m_matrix[10][23] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\m_blake2.m_hash256.v_q[4][2] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\m_blake2.m_hash256.m_matrix[6][8] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\m_blake2.m_hash256.v_q[10][27] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(\m_io.m_config.ll_q[22] ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\m_blake2.m_hash256.v_q[13][1] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\m_blake2.m_hash256.m_matrix[1][31] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\m_blake2.m_hash256.m_matrix[6][23] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\m_blake2.m_hash256.v_q[12][31] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[10] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\m_io.m_config.kk_q[2] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\m_blake2.m_hash256.v_q[9][9] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\m_blake2.m_hash256.m_matrix[5][25] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\m_blake2.m_hash256.m_matrix[5][25]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\m_blake2.m_hash256.m_matrix[13][28] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\m_blake2.m_hash256.m_matrix[11][8] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\m_blake2.m_hash256.m_matrix[2][7] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\m_blake2.m_hash256.m_matrix[4][3] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[50] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[55] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\m_blake2.m_hash256.m_matrix[11][16] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\m_io.m_config.ll_q[8] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(\m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\m_blake2.m_hash256.m_matrix[2][6] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[34] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\m_blake2.m_hash256.block_idx_plus_one_q[6] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(\m_blake2.m_hash256.v_q[13][12] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\m_blake2.m_hash256.h_flat[125] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(\m_blake2.m_hash256.m_matrix[1][3] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\m_blake2.m_hash256.v_q[11][18] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(\m_blake2.m_hash256.m_matrix[8][4] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\m_blake2.m_hash256.v_q[10][26] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\m_blake2.m_hash256.slow_output_q ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\m_blake2.m_hash256.m_matrix[5][16] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\m_blake2.m_hash256.m_matrix[2][28] ),
    .X(net1905));
 sky130_fd_sc_hd__buf_1 fanout1 (.A(\m_io.en_q ),
    .X(net1906));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_A (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(ena));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_A1 (.DIODE(\hash[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[0]_sky130_fd_sc_hd__or2_2_B_B  (.DIODE(\hash[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\hash[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[0]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\hash[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D_sky130_fd_sc_hd__a22o_2_X_B2 (.DIODE(\hash[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[3]_sky130_fd_sc_hd__mux2_1_A0_A0  (.DIODE(\hash[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\hash[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\hash[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[11]_sky130_fd_sc_hd__o22a_2_A2_X  (.DIODE(\hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\hash[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2_A1  (.DIODE(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[3]_sky130_fd_sc_hd__mux2_1_A0_X  (.DIODE(\hash[3]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D_sky130_fd_sc_hd__a22o_2_X_B2 (.DIODE(\hash[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__mux2_1_A0_A0  (.DIODE(\hash[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\hash[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\hash[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__o22a_2_A2_X  (.DIODE(\hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\hash[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2_A1  (.DIODE(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_B  (.DIODE(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__mux2_1_A0_X  (.DIODE(\hash[4]_sky130_fd_sc_hd__mux2_1_A0_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_B2 (.DIODE(\hash[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[5]_sky130_fd_sc_hd__mux2_1_A1_A1  (.DIODE(\hash[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\hash[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\hash[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[13]_sky130_fd_sc_hd__o22a_2_A2_X  (.DIODE(\hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__a21bo_2_A2_A1  (.DIODE(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[5]_sky130_fd_sc_hd__mux2_1_A1_X  (.DIODE(\hash[5]_sky130_fd_sc_hd__mux2_1_A1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D_sky130_fd_sc_hd__a22o_2_X_B2 (.DIODE(\hash[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[6]_sky130_fd_sc_hd__or2_2_B_B  (.DIODE(\hash[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\hash[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\hash[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_B2 (.DIODE(\hash[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\hash[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\hash[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[7]_sky130_fd_sc_hd__and2_2_B_B  (.DIODE(\hash[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_B_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_A  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2_sky130_fd_sc_hd__nor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X_C  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[16]_sky130_fd_sc_hd__and4_2_C_D  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_C_sky130_fd_sc_hd__a21o_2_X_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__and4_2_C_C  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[7]_sky130_fd_sc_hd__a22o_2_B2_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__and4_2_B_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__a221o_2_A1_B2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__and3_2_B_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[27]_sky130_fd_sc_hd__a31o_2_B1_B1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[34]_sky130_fd_sc_hd__a22oi_2_B2_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[30]_sky130_fd_sc_hd__a31o_2_B1_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[28]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__a31o_2_B1_A3  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__and2_2_A_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[33]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[39]_sky130_fd_sc_hd__a31o_2_B1_A3  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[37]_sky130_fd_sc_hd__and2_2_A_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__a31o_2_B1_A3  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__and2_2_A_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[42]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[48]_sky130_fd_sc_hd__a31o_2_B1_A3  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[46]_sky130_fd_sc_hd__and2_2_A_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_A_N  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__o21ai_2_A1_A2_sky130_fd_sc_hd__and3_2_X_C  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[7]_sky130_fd_sc_hd__and4_2_C_D  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_A2  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__and2_2_X_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[57]_sky130_fd_sc_hd__a221o_2_B2_A1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[51] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[51] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__and3_2_B_B  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[51] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[51]_sky130_fd_sc_hd__a31o_2_B1_B1  (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[51] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C  (.DIODE(\m_blake2.m_hash256.f_finished ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a31o_2_X_B1_sky130_fd_sc_hd__and3b_2_X_A_N  (.DIODE(\m_blake2.m_hash256.f_finished ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.f_finished_sky130_fd_sc_hd__and2_2_X_X  (.DIODE(\m_blake2.m_hash256.f_finished ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.f_finished_q_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.f_finished ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A2_sky130_fd_sc_hd__nor2_2_Y_B  (.DIODE(\m_blake2.m_hash256.f_finished ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout500_A (.DIODE(\m_blake2.m_hash256.first_block_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout494_A (.DIODE(\m_blake2.m_hash256.first_block_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout489_A (.DIODE(\m_blake2.m_hash256.first_block_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout486_A (.DIODE(\m_blake2.m_hash256.first_block_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.first_block_q_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.first_block_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_A (.DIODE(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[44]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[1]_sky130_fd_sc_hd__o21a_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X  (.DIODE(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_block_last_sky130_fd_sc_hd__a22o_2_B2_B1_sky130_fd_sc_hd__nor2_2_Y_A (.DIODE(\m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_A (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout305_A (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout304_A (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout480_A (.DIODE(\m_blake2.m_hash256.fsm_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout479_A (.DIODE(\m_blake2.m_hash256.fsm_q[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_A (.DIODE(\m_blake2.m_hash256.fsm_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(\m_blake2.m_hash256.fsm_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.fsm_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y  (.DIODE(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[14] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y  (.DIODE(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_A1  (.DIODE(\m_blake2.m_hash256.g_b[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1_A2  (.DIODE(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B  (.DIODE(\m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_B2  (.DIODE(\m_blake2.m_hash256.g_b[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A  (.DIODE(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1  (.DIODE(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X  (.DIODE(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_B  (.DIODE(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2  (.DIODE(\m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_Y  (.DIODE(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y  (.DIODE(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B  (.DIODE(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_Y  (.DIODE(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[25]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nand2b_2_Y_B  (.DIODE(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__xnor2_2_B_A  (.DIODE(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N  (.DIODE(\m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_X_A  (.DIODE(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1  (.DIODE(\m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A  (.DIODE(\m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_b[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_b[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.g_b[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__and2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_Y  (.DIODE(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_X  (.DIODE(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[11]_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(\m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[7]_sky130_fd_sc_hd__a21o_2_X_A1  (.DIODE(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[6]_sky130_fd_sc_hd__a211o_2_X_A1  (.DIODE(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1_sky130_fd_sc_hd__nor2_2_Y_Y  (.DIODE(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1  (.DIODE(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[2]_sky130_fd_sc_hd__a211o_2_X_A1  (.DIODE(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[0]_sky130_fd_sc_hd__a211o_2_X_A1  (.DIODE(\m_blake2.m_hash256.g_c_buf[3]_sky130_fd_sc_hd__a21o_2_X_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_d[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_X  (.DIODE(\m_blake2.m_hash256.g_d[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D  (.DIODE(\m_blake2.m_hash256.g_d[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_X  (.DIODE(\m_blake2.m_hash256.g_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(\m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(\m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X  (.DIODE(\m_blake2.m_hash256.g_idx_next[0]_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X  (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3_2_A_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X  (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__and3b_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y  (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X  (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout412_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_A (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X  (.DIODE(\m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__or3b_2_A_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X  (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__and2b_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y  (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y  (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y  (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y  (.DIODE(\m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y  (.DIODE(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_A (.DIODE(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.h_flat[131] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__mux2_1_A0_A0  (.DIODE(\m_blake2.m_hash256.h_flat[131] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.h_flat[131] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[131] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.h_flat[132] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__mux2_1_A0_A0  (.DIODE(\m_blake2.m_hash256.h_flat[132] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.h_flat[132] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[132]_sky130_fd_sc_hd__a22o_2_A1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[132] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.h_flat[133] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__mux2_1_A0_A0  (.DIODE(\m_blake2.m_hash256.h_flat[133] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.h_flat[133] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__a22o_2_A1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[133] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.h_flat[134] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__mux2_1_A0_A0  (.DIODE(\m_blake2.m_hash256.h_flat[134] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.h_flat[134] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__a22o_2_A1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[134] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand2_2_B_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[247]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[239]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_A1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o32a_2_X_B2  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_A1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_2_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[107]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_A  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_B2  (.DIODE(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2_sky130_fd_sc_hd__nand2_2_Y_Y  (.DIODE(\m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_B2  (.DIODE(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_B2  (.DIODE(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_Y  (.DIODE(\m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_A1  (.DIODE(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_A1  (.DIODE(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y_Y  (.DIODE(\m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_A (.DIODE(\m_blake2.m_hash256.last_block_q ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(\m_blake2.m_hash256.last_block_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[42]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(\m_blake2.m_hash256.last_block_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.last_block_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.last_block_q_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.last_block_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_X  (.DIODE(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2  (.DIODE(\m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X_sky130_fd_sc_hd__xnor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(\m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__inv_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[13]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[30]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_A2_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[31]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[14]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.a_q[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[15]_sky130_fd_sc_hd__a21oi_2_A1_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_A_sky130_fd_sc_hd__a21bo_2_X_A1_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[16]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.a_q[18]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__a21o_2_A1_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[6]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[22]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.a_q[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[23]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.a_q[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and3_2_C_C  (.DIODE(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__a21o_2_B1_B1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__nand2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[14]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X  (.DIODE(\m_blake2.m_hash256.m_g.a_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__a21boi_2_A1_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[23]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X  (.DIODE(\m_blake2.m_hash256.m_g.a_q[6]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor3b_2_C_N_Y_sky130_fd_sc_hd__o21ba_2_A1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21oi_2_A2_Y_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[26]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X  (.DIODE(\m_blake2.m_hash256.m_g.a_q[9]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__o31a_2_B1_X_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][10]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][12]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_C  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_A2  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand3_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][15]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][17]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][16]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__and2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][18]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][19]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__and2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[18]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__and2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][23]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][23]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][22]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[22]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][25]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][27]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[7]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[22]_sky130_fd_sc_hd__nand2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2_sky130_fd_sc_hd__o21bai_2_Y_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_A2  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A3_sky130_fd_sc_hd__a21o_2_X_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_C  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_A2  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__a21bo_2_B1_N_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[31]_sky130_fd_sc_hd__nand3b_2_A_N_Y_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][7]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a21o_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.b_q[6]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[21]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][3]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.c_q[0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__a41o_2_A2_X_sky130_fd_sc_hd__a21bo_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[16]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.c_q[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__o211a_2_A1_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.c_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[19]_sky130_fd_sc_hd__a221o_2_A1_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.c_q[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__o211a_2_A1_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[7]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__o211a_2_C1_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B_sky130_fd_sc_hd__o21a_2_X_A1  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_B_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[4]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2b_2_X_A_N_sky130_fd_sc_hd__nor2_2_Y_A  (.DIODE(\m_blake2.m_hash256.m_g.c_q[3]_sky130_fd_sc_hd__a221oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][19]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nand2b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[19]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__and2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.m_g.d_q[11]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][20]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][20]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][20]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[12]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][23]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][23]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][23]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[23]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_A1_A2  (.DIODE(\m_blake2.m_hash256.m_g.d_q[15]_sky130_fd_sc_hd__xnor2_2_B_Y_sky130_fd_sc_hd__xnor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[24]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[16]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][25]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][25]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__nand2b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[25]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_A_N  (.DIODE(\m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.c_q[17]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a21oi_2_B1_A2  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__and2_2_X_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[11]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__a21oi_2_B1_Y_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__nor2_2_Y_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[20]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[30]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__a32o_2_B2_A1_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[28]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__xnor2_2_Y_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[21]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[17]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.d_q[9]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[0]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[10]_sky130_fd_sc_hd__and2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[11]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[12]_sky130_fd_sc_hd__and2b_2_A_N_A_N  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[12] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__inv_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[13]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[13] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[14]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[15]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[15] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[16]_sky130_fd_sc_hd__and2b_2_A_N_A_N  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[16] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xnor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[17]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__inv_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[18]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[18] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__nand3b_2_A_N_A_N  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[19]_sky130_fd_sc_hd__a21bo_2_B1_N_B1_N  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[19] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__and3_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21oi_2_B1_B1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[1]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[20]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[21]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[21] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[23]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[23] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[29]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__o21bai_2_B1_N_Y_sky130_fd_sc_hd__o311a_2_C1_A1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__nand3_2_C_Y_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__xor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_Y_sky130_fd_sc_hd__o311a_2_B1_A1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[28]_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a21o_2_B1_X_sky130_fd_sc_hd__o211ai_2_C1_A1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__a21oi_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_Y_sky130_fd_sc_hd__a21boi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[24]_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nand3_2_A_Y_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__xnor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[25]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[26]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[26] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[27]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[27] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[28]_sky130_fd_sc_hd__and2b_2_A_N_A_N  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[28] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[29]_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[29] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[30]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[31]_sky130_fd_sc_hd__xor2_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[31] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[31]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[31] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__and3_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[3]_sky130_fd_sc_hd__a21oi_2_B1_B1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[4]_sky130_fd_sc_hd__and2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__inv_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[5]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[6]_sky130_fd_sc_hd__and2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__and3_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[7]_sky130_fd_sc_hd__a21oi_2_B1_B1  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__nand2b_2_B_B  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[8]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.m_add_1.x2_i[9]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_blake2.m_hash256.m_g.m_add_1.x2_i[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X_sky130_fd_sc_hd__and3_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X  (.DIODE(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(\m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__and2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X  (.DIODE(\m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X_sky130_fd_sc_hd__inv_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X  (.DIODE(\m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X  (.DIODE(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a22o_2_B2_A1  (.DIODE(\m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y  (.DIODE(\m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__nand2b_2_A_N_A_N  (.DIODE(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y  (.DIODE(\m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X  (.DIODE(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N  (.DIODE(\m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_A  (.DIODE(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_A_N  (.DIODE(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y  (.DIODE(\m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_A (.DIODE(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_A (.DIODE(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y  (.DIODE(\m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__nand2b_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout83_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout75_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_X_sky130_fd_sc_hd__or4_2_B_X_sky130_fd_sc_hd__o22a_2_B1_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o31a_2_A1_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_B1_sky130_fd_sc_hd__or2_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_5_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_D_6_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_1_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_2_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X  (.DIODE(\m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o41a_2_A3_X_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__and4_2_D_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X  (.DIODE(\m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_X_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X  (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_3_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X  (.DIODE(\m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__nor3_2_C_Y_sky130_fd_sc_hd__and4_2_C_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y  (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_A_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout39_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout37_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y  (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_B_Y_sky130_fd_sc_hd__nor2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_A (.DIODE(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout317_A (.DIODE(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_A (.DIODE(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y  (.DIODE(\m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__nand2b_2_A_N_A_N  (.DIODE(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y  (.DIODE(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__nand2b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_Y_sky130_fd_sc_hd__xor2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X_sky130_fd_sc_hd__and2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X  (.DIODE(\m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A_sky130_fd_sc_hd__or2_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1_A1  (.DIODE(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__a21oi_2_B1_A2  (.DIODE(\m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X  (.DIODE(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_C  (.DIODE(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X  (.DIODE(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B  (.DIODE(\m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X  (.DIODE(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__o211ai_2_A2_C1  (.DIODE(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2  (.DIODE(\m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X_sky130_fd_sc_hd__xnor2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X  (.DIODE(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B1  (.DIODE(\m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X  (.DIODE(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_Y_sky130_fd_sc_hd__and2b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(\m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__mux4_2_A0_S1  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__xor2_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1_B  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_C  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__o211a_2_C1_B1  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_C  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_C  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[23]_sky130_fd_sc_hd__o311a_2_X_A3  (.DIODE(\m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A1  (.DIODE(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[8]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_B_X_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__xor2_2_B_X  (.DIODE(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[20]_sky130_fd_sc_hd__xnor2_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_A1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__o22a_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2_sky130_fd_sc_hd__or2_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__o22a_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__o22a_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[10]_sky130_fd_sc_hd__xnor2_2_A_B_sky130_fd_sc_hd__and2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][12]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[4]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_B  (.DIODE(\m_blake2.m_hash256.v_q[12][12]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][13]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][13]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][13]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[5]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__or4_2_A_B_sky130_fd_sc_hd__xor2_2_X_B  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_X_sky130_fd_sc_hd__o21ai_2_A2_B1_sky130_fd_sc_hd__nand2b_2_Y_A_N  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__and2b_2_A_N_X_sky130_fd_sc_hd__a31o_2_B1_A3  (.DIODE(\m_blake2.m_hash256.v_q[12][13]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][15]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][15]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][15]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[7]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__xor2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[15]_sky130_fd_sc_hd__nand3_2_A_B_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(\m_blake2.m_hash256.v_q[12][15]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][21]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[13]_sky130_fd_sc_hd__xor2_2_B_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][5]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][5]_sky130_fd_sc_hd__mux2_1_A0_A1  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][5]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[29]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__xor2_2_A_X  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__xnor2_2_A_B  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o21ai_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[5]_sky130_fd_sc_hd__xor2_2_A_B_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__a21o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[12][5]_sky130_fd_sc_hd__mux2_1_A1_A0 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][20]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][29]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1_sky130_fd_sc_hd__nor2_2_Y_Y  (.DIODE(\m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(\m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nand3_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B  (.DIODE(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_B  (.DIODE(\m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_X_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[4]_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2_sky130_fd_sc_hd__and2_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_A (.DIODE(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[0]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__o31a_2_A2_B1  (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__or2_2_X_X  (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__a32o_2_A1_B1  (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y  (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y  (.DIODE(\m_io.m_config.cfg_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__or2_2_X_B_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_7_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2 (.DIODE(\m_io.m_config.data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[0]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_6_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2 (.DIODE(\m_io.m_config.data_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[57]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[1]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_5_D_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2 (.DIODE(\m_io.m_config.data_i[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[58]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[2]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_4_D_sky130_fd_sc_hd__a22o_2_X_A1 (.DIODE(\m_io.m_config.data_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[3]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_3_D_sky130_fd_sc_hd__a22o_2_X_A1 (.DIODE(\m_io.m_config.data_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[4]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_2_D_sky130_fd_sc_hd__o22a_2_X_A1 (.DIODE(\m_io.m_config.data_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[5]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_1_D_sky130_fd_sc_hd__a22o_2_X_A1 (.DIODE(\m_io.m_config.data_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[62]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[6]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_uo_out_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a22o_2_X_A1 (.DIODE(\m_io.m_config.data_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.data_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.data_i[7]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.data_i[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_data[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_A0  (.DIODE(\m_io.m_config.data_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X  (.DIODE(\m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__and3_2_B_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[3]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_io.m_config.kk_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_A1  (.DIODE(\m_io.m_config.kk_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.kk_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[4]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_io.m_config.kk_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1_A1  (.DIODE(\m_io.m_config.kk_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.kk_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nand2_2_A_A  (.DIODE(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_A0  (.DIODE(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_A (.DIODE(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1_sky130_fd_sc_hd__nand2_2_Y_Y  (.DIODE(\m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[60]_sky130_fd_sc_hd__a211o_2_A1_C1  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[56]_sky130_fd_sc_hd__a211o_2_A1_C1  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_Y  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X  (.DIODE(\m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_C1_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__or2_2_A_X ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[56]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_io.m_config.ll_q[56] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.ll_q[56] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[56]_sky130_fd_sc_hd__a211o_2_A1_A1  (.DIODE(\m_io.m_config.ll_q[56] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[48]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.ll_q[56] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[59]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_io.m_config.ll_q[59] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[59]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.ll_q[59] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[59]_sky130_fd_sc_hd__a221o_2_B2_B2  (.DIODE(\m_io.m_config.ll_q[59] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[51]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.ll_q[59] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[63]_sky130_fd_sc_hd__or2_2_A_A  (.DIODE(\m_io.m_config.ll_q[63] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[63]_sky130_fd_sc_hd__dfxtp_2_Q_Q  (.DIODE(\m_io.m_config.ll_q[63] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[63]_sky130_fd_sc_hd__a22oi_2_B2_B2  (.DIODE(\m_io.m_config.ll_q[63] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A1  (.DIODE(\m_io.m_config.ll_q[63] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y  (.DIODE(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__xor2_2_A_X_sky130_fd_sc_hd__a21oi_2_B1_A1  (.DIODE(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[0]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(\m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y  (.DIODE(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_B1_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[5]_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(\m_io.m_config.nn_q[5]_sky130_fd_sc_hd__inv_2_A_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(rst_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(ui_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(ui_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(ui_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(ui_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(ui_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(ui_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(ui_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(ui_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(uio_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(uio_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(uio_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(uio_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(uio_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout615_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_X (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout16_X (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_X (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_X (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_X (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_X (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_X (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_X (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[2]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout24_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_X (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_X (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_X (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_X (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_X (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_X (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[23]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_X (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_X (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout46_X (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_X (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_X (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_X (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout56_X (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_X (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_X (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_X (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[27]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[18]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_X (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_X (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_X (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_X (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[30]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_X (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[11]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_X (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[15]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_X (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[26]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_X (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[22]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[14]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[4]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[28]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[12]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[20]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[29]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[21]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[13]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_X (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[3]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[19]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[0]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[8]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[24]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[16]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[9]_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[25]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[17]_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_y_buf[1]_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_X (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_X (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_X (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_X (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_X (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_X (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_X (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_X (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_B1  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_A2  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_B1  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_A2  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_X (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_B1  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_A_sky130_fd_sc_hd__or2_2_X_B  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][0]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_X (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_B1  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_X (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_A  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_D1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_X (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_X (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_X (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_X (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_X (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_B1  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_X (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X_A2  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_X (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][7]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_X (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_X (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A3_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_X (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_X (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_X (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_X (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__a22oi_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][6]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_X (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_X (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_X (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_X (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a21o_2_X_A2  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_X (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_X (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A3_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_X (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B1_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A1_sky130_fd_sc_hd__a221oi_2_Y_B1  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_X (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A1_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A2  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_X (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__a22o_2_B2_A1_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][4]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_X_sky130_fd_sc_hd__o21a_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__a32o_2_X_A2_sky130_fd_sc_hd__a2111oi_2_Y_A2  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][5]_sky130_fd_sc_hd__o22ai_2_A1_B2_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_X (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__a21oi_2_A1_B1_sky130_fd_sc_hd__and3_2_X_B_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__and3_2_C_B_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[0]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ba_2_X_A2_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32ai_2_Y_A2_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][1]_sky130_fd_sc_hd__o32a_2_B2_A2_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o2bb2a_2_B2_A1_N_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__nor3_2_Y_C_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_X (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a0[28]_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__o32a_2_X_A1_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][3]_sky130_fd_sc_hd__o22a_2_A1_B2_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__a22o_2_X_B1  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_X_sky130_fd_sc_hd__or2_2_B_A_sky130_fd_sc_hd__o32a_2_X_A3_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_C1_A2_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_X (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_X (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][20]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_X (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_X (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][31]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_X (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_X (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_X (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][31]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_X (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_X (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[33]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_X (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[37]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_A2  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_X (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__a32o_2_A1_B1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_X (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__a32o_2_A1_B1  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_X (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__a221o_2_A1_B2  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__a32o_2_A1_B1  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_B1  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__a221o_2_A1_B2  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__a32o_2_A1_B1  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_X (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][23]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][15]_sky130_fd_sc_hd__o22a_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][29]_sky130_fd_sc_hd__o22a_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][22]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][14]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_X (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_B2  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__o22a_2_A1_B1  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_X (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[11]_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[22]_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[12]_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[8]_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[26]_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[18]_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[17]_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_X (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[19]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[15]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[14]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[5]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[13]_sky130_fd_sc_hd__o32a_2_X_B1  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[9]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[1]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[10]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[16]_sky130_fd_sc_hd__o22a_2_X_A2  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_X (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_B1_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B2_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_X (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_C1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_X (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_C1  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1_C1  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_X (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_C1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][21]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21o_2_X_B1_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][15]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_X (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][23]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a211o_2_A2_C1  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_X (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[26]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[10]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[25]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_X (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[13]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[21]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[15]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[31]_sky130_fd_sc_hd__o21a_2_X_A1  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[23]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_X (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_B2_sky130_fd_sc_hd__a21o_2_X_B1  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_X (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout183_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[27]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[11]_sky130_fd_sc_hd__inv_2_Y_A_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_X (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_D_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__a221o_2_A1_B2  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__a221o_2_A1_B2  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_A_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_X (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][12]_sky130_fd_sc_hd__a221o_2_A1_B2  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[7]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_B1_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_X (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_X_sky130_fd_sc_hd__a221o_2_B1_B2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_A1_N  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_A1_N  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_X (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[173]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_A1_N  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[15]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][27]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_B_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][24]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_X (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_B_sky130_fd_sc_hd__o21a_2_X_B1  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[30]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_X (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][2]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][10]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][17]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][1]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][25]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][9]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_X (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[251]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][8]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][19]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][18]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_X (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][26]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_X (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][22]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][4]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][28]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][24]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][14]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][3]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_X (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][13]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][5]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][20]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_B1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][30]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][12]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_X (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][19]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][17]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][26]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][10]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][25]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][29]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][31]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][23]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][13]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][15]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][20]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][30]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][22]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][21]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][12]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][24]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][28]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][14]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_X (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][11]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][27]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][18]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][25]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][9]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][17]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][2]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][1]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][0]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_X (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][29]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][12]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][3]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][24]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][4]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][28]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][14]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][6]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][27]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][16]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][18]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_X (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][0]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][2]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][1]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][9]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_X (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][6]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][4]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][3]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][16]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][27]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][11]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_X (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][19]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][17]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][20]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][22]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][14]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][24]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][28]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_X (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][30]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][12]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][29]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][18]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][26]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][18]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][10]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][16]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][25]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][17]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][8]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][0]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][24]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][20]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][12]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][2]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_X (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][19]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][3]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][11]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][4]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][28]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][21]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_X (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][26]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][18]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][10]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][16]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][17]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_X (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][12]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][24]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_X (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][22]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][14]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][15]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][29]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][30]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][23]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_X (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][27]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][19]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][11]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][31]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][28]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][13]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][21]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_X (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][0]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][17]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][25]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][2]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][26]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][9]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][1]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_X (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][31]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][3]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][4]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][28]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][6]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][14]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_X (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_X (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][13]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][12]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][22]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][20]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][31]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][23]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][15]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][1]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][16]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][8]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][0]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][20]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][12]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][2]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_X (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][31]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][22]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][23]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][6]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][15]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][27]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][7]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][3]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][4]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][13]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_X (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_B1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[10]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_C1_sky130_fd_sc_hd__o211a_2_X_B1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[0]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_X (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[29]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A1_sky130_fd_sc_hd__o211a_2_X_B1  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_C_sky130_fd_sc_hd__o211a_2_X_B1  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout240_X (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[9]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_D1_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[17]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o221a_2_X_B1  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_X (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[8]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[51]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[41]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_X (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[37]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[60]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[14]_sky130_fd_sc_hd__or2_2_A_B  (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_X (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__a311o_2_A1_A3  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__a311o_2_A1_A3  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][11]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_B  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__o31a_2_A1_A3  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_B  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][25]_sky130_fd_sc_hd__a22o_2_A1_B2  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__a32o_2_A1_A3  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_X (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][16]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__a32o_2_A1_A3  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][2]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][26]_sky130_fd_sc_hd__a32o_2_A1_A3  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][18]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][10]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][17]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][0]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][9]_sky130_fd_sc_hd__a221o_2_A1_B2  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_X (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][6]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][30]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][29]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][22]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][3]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][15]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[21]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[28]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][13]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__a32o_2_A1_A3  (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_X (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][7]_sky130_fd_sc_hd__a22o_2_A1_B2  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[31]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__a32o_2_A1_A3  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[24]_sky130_fd_sc_hd__a221o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_X (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][13]_sky130_fd_sc_hd__o22a_2_A1_B2  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout253_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[19]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_A2_sky130_fd_sc_hd__or2_2_X_B  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[16]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][2]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][0]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][1]_sky130_fd_sc_hd__o22a_2_A1_B2  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[9]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[10]_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_X (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[19]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[24]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[2]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_A1  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_X (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[18]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][27]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_A1  (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_X (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[223]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[7]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[5]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][13]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a221o_2_A2_A1  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[20]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_X (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][31]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[12]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[3]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_A1  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[6]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[14]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_B2  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[28]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_X (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][19]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[59]_sky130_fd_sc_hd__a221o_2_B2_A2  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][26]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][10]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[26]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_A2  (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_X (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[43]_sky130_fd_sc_hd__a221o_2_B2_A2  (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[16]_sky130_fd_sc_hd__a22o_2_B2_A2  (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[48]_sky130_fd_sc_hd__a22oi_2_B2_A2  (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_X (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_B2  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_A1  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[92]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_A1  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_B2  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_B2  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_X (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[61]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211a_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[47]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[43]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__o221a_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[49]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o211ai_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_B2  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_A1  (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_X (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][8]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[27]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[25]_sky130_fd_sc_hd__a221o_2_B2_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[25]_sky130_fd_sc_hd__a21oi_2_Y_A2_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[26]_sky130_fd_sc_hd__a221o_2_B2_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][10]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_X (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][29]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_B1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[15]_sky130_fd_sc_hd__a221o_2_B2_C1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][21]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][23]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[20]_sky130_fd_sc_hd__a221o_2_B2_C1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][22]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_A  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__and4_2_X_A  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_X (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[8]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[19]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[24]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[3]_sky130_fd_sc_hd__or4_2_X_A_sky130_fd_sc_hd__o221a_2_X_C1  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__a221o_2_A1_C1  (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_X (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[5]_sky130_fd_sc_hd__a211o_2_X_C1_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[21]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[23]_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[12]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[28]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[4]_sky130_fd_sc_hd__or3_2_X_C_sky130_fd_sc_hd__a22o_2_X_B2  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[14]_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[6]_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_B1_sky130_fd_sc_hd__a221o_2_X_C1  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_X (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[29]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o32a_2_X_A3  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[30]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[4]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A3  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[1]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B2  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_B2  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a2bb2o_2_B1_A1_N  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o22a_2_X_B2  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[0]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A2_N_sky130_fd_sc_hd__o2bb2a_2_X_B1  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_X (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[31]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[13]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[2]_sky130_fd_sc_hd__a2111o_2_X_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[1]_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[18]_sky130_fd_sc_hd__o2bb2a_2_X_B1_sky130_fd_sc_hd__a221o_2_X_A2  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_X (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_A1  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_B2  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_X (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__a21oi_2_A1_A2  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_B2  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_A1  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_X (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__a21oi_2_A1_A2  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_X (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_B2  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_A1  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__a211oi_2_A1_A2  (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_X (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3_2_X_C_sky130_fd_sc_hd__a21o_2_X_A1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__a211oi_2_A1_A2  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_X (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_A1  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21bo_2_A2_A1  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[2]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2_B2  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_X (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[39]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_A1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_X (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[83]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[99]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[91]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[95]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_X (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_B2  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__a211oi_2_A1_A2  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_A1  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_A1  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_A1  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_X (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[90]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_X (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21boi_2_A2_A1  (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_A1  (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_X (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_X (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_X (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_A1  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[53]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_X (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][8]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][0]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][9]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][2]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][1]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_X (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][4]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][6]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][3]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_X (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][16]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_X (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][20]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][12]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_A1  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_1_A  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_X (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][27]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][22]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][15]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][23]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_X (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][11]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][31]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][13]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout307_X (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[20]_sky130_fd_sc_hd__a221o_2_B2_B1  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[22]_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_A2  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[45]_sky130_fd_sc_hd__a22oi_2_B2_B1  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[56]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[60]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[46]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[4]_sky130_fd_sc_hd__o2bb2a_2_A1_N_A2_N  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[35]_sky130_fd_sc_hd__a22oi_2_B2_B1  (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout314_X (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout313_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout310_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_X (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[60]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[12]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_X (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[195]_sky130_fd_sc_hd__a21o_2_A1_A2  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[227]_sky130_fd_sc_hd__a21o_2_A1_A2  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[163]_sky130_fd_sc_hd__a21o_2_A1_A2  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[208]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_X (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[164]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[230]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[182]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_X (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1_A2  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout327_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_X (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout334_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[75]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[115]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[15]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[19]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_X (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout340_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout342_X (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout332_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout326_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout346_X (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout345_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[106]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a31o_2_A3_B1  (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][8]_sky130_fd_sc_hd__a32o_2_A1_A2  (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_B1_X_sky130_fd_sc_hd__or3_2_C_A  (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_C1  (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_B1  (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][1]_sky130_fd_sc_hd__a32o_2_A1_A2  (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_C1  (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_X (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][27]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][11]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[16]_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a211o_2_X_A2  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[16]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__and2_2_X_A  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][8]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A2_sky130_fd_sc_hd__a21o_2_X_A1  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[8]_sky130_fd_sc_hd__o22a_2_X_A1_sky130_fd_sc_hd__a2bb2o_2_X_A1_N  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][24]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(net349));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout350_X (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][27]_sky130_fd_sc_hd__a22o_2_A1_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][11]_sky130_fd_sc_hd__a221o_2_A1_A2  (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout349_A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a211o_2_A2_C1  (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_B1  (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_C1  (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][12]_sky130_fd_sc_hd__a32o_2_A1_A2  (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_X (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout353_A (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][4]_sky130_fd_sc_hd__a32o_2_A1_A2  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_A1  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21oi_2_A2_B1  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[77]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_A2_C1  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_C1  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[85]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a211oi_2_A2_C1  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[20]_sky130_fd_sc_hd__and2_2_X_A  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][14]_sky130_fd_sc_hd__a311o_2_A1_A2  (.DIODE(net354));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_X (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[71]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a21o_2_A2_B1  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_X_sky130_fd_sc_hd__a221o_2_B1_C1  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_B  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[30]_sky130_fd_sc_hd__a22o_2_X_A1  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_B  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__nand2_2_A_Y_sky130_fd_sc_hd__a31o_2_A2_A1  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][25]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][3]_sky130_fd_sc_hd__a22o_2_A1_A2_sky130_fd_sc_hd__and2_2_X_A  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[23]_sky130_fd_sc_hd__o311a_2_X_C1  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][19]_sky130_fd_sc_hd__a311o_2_A1_A2  (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_X (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_X (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_b[17]_sky130_fd_sc_hd__o22a_2_X_B1_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][1]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout370_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout365_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__a211oi_2_A1_C1  (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_X (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[13][11]_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[15][11]_sky130_fd_sc_hd__o21ai_2_A1_A2  (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_d[11]_sky130_fd_sc_hd__a21oi_2_Y_A1_sky130_fd_sc_hd__o21ai_2_Y_A2  (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][11]_sky130_fd_sc_hd__mux2_1_A0_1_S  (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout376_A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_X (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__o31a_2_A1_A2  (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][5]_sky130_fd_sc_hd__o21a_2_A1_A2  (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_X (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout397_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout399_X (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__a211o_2_A1_C1  (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_X (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[79]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_A2_B2  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[70]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[78]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_B2  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[81]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_B2  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[41]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_A1  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o221a_2_B1_A1  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22ai_2_A2_B2  (.DIODE(net400));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_X (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__or3_2_B_A_sky130_fd_sc_hd__o211a_2_X_B1  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_D_X_sky130_fd_sc_hd__or4_2_D_C_sky130_fd_sc_hd__a32o_2_X_B2  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__or4_2_C_D_sky130_fd_sc_hd__o311a_2_X_B1  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[5]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__a311o_2_B1_A2  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__or3_2_B_X_sky130_fd_sc_hd__o211a_2_A2_C1  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[1]_sky130_fd_sc_hd__o311a_2_A1_B1  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__o31a_2_A1_X_sky130_fd_sc_hd__nor4_2_B_D_sky130_fd_sc_hd__o311a_2_X_B1  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[2]_sky130_fd_sc_hd__mux2_1_A1_X_sky130_fd_sc_hd__a221oi_2_A2_A1  (.DIODE(net401));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_X (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[0]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__a211o_2_A1_A2  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__a211oi_2_A1_A2  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[1]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net402));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_X (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_A1  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout401_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__a221o_2_A1_B1  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_X (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__o2bb2a_2_A2_N_A1_N  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22oi_2_A2_A1  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_A2_A1  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a21o_2_A2_A1  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_X (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[1][4]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a22o_2_B1_B2  (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__a22o_2_A1_B1  (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[45]_sky130_fd_sc_hd__or2_2_B_X_sky130_fd_sc_hd__a22o_2_A2_B2  (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A0_X_sky130_fd_sc_hd__a2bb2o_2_B1_B2  (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout407_X (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][14]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][25]_sky130_fd_sc_hd__or3_2_B_A  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_1_A  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[9]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__a22o_2_A2_B1_sky130_fd_sc_hd__or3_2_X_A  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[7]_sky130_fd_sc_hd__or4_2_A_1_X_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.round_q[0]_sky130_fd_sc_hd__or3_2_C_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nor3_2_B_C_sky130_fd_sc_hd__o31a_2_X_A1  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_B  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][9]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y_B  (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_X (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][11]_sky130_fd_sc_hd__nand2_2_A_B_sky130_fd_sc_hd__and3_2_X_A  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[11][27]_sky130_fd_sc_hd__a22o_2_A1_B2  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][23]_sky130_fd_sc_hd__a22o_2_B1_A1  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][27]_sky130_fd_sc_hd__o31a_2_A2_A1  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_A  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][19]_sky130_fd_sc_hd__o21a_2_A1_B1  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][5]_sky130_fd_sc_hd__o31a_2_A1_B1  (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_X (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][18]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][10]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_A1_B1_N  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][16]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][25]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][17]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout410_X (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][20]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][24]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][12]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][26]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_X (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][11]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][29]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][30]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][23]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][22]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][15]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][14]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout412_X (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][31]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][19]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][27]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][28]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][13]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][21]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[0][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_X (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__and2_2_A_X_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_1_A1  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][16]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_X (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][20]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][12]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout413_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_X (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][11]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][22]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][15]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][23]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_X (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][27]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][31]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][13]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[2][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_X (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][26]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][18]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][10]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][16]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][8]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][25]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][17]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout418_X (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][20]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][12]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][24]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__o21ai_2_B1_Y_sky130_fd_sc_hd__o21ai_2_B1_1_A1  (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__a21bo_2_B1_N_X_sky130_fd_sc_hd__o21ai_2_B1_A1  (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__o21a_2_A1_X_sky130_fd_sc_hd__o21ba_2_B1_N_A1  (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout417_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_X (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][27]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][29]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][7]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][30]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][15]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][14]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][6]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][23]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][22]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout420_X (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][11]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][19]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][31]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout419_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][28]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][21]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__mux2_1_X_S  (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_X (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[38]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[32]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[57]_sky130_fd_sc_hd__a21oi_2_A1_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[29]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[20]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[53]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout422_X (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[47]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout421_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[35]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[11]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__a21oi_2_Y_B1  (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_X (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[55]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[21]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[19]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[43]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[45]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[36]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and3b_2_X_B  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[13]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[34]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout427_X (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[56]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout425_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout424_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout426_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.ready_v_o_sky130_fd_sc_hd__o21a_2_X_B1_sky130_fd_sc_hd__mux2_1_A1_A0  (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[4]_sky130_fd_sc_hd__o21ai_2_A1_B1  (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.block_idx_plus_one_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_B_sky130_fd_sc_hd__o21ai_2_Y_B1  (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_X (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[89]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[121]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[40]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[64]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[96]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[26]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[33]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout428_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_X (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[194]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[153]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[177]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[2]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[2]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[1]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[169]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[233]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[241]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_X (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[225]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[202]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[161]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout430_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout429_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_X (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[211]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[226]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[154]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[242]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[210]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[186]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_X (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout432_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout433_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[88]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[44]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[84]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[52]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[116]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[20]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_X (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[166]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[198]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[148]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[36]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[124]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[37]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[117]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[5]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[21]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[28]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_X (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[67]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[94]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[62]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[46]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[119]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[55]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[87]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[102]_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[126]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[38]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_X (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout439_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout440_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[180]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[172]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[190]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[222]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[212]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[244]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[214]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_X (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[221]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout441_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[7]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[22]_sky130_fd_sc_hd__and2_2_B_A  (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout438_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout437_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout443_X (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout436_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout435_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout442_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout431_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout434_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_X (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[138]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[232]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_B1_sky130_fd_sc_hd__a21oi_2_Y_A1  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21ai_2_Y_A1  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__a21oi_2_B1_A1  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__xor2_2_B_A  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_A1  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_X (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[236]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout448_X (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout447_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[170]_sky130_fd_sc_hd__and3_2_C_A  (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout446_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_X (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[58]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[49]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[41]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[18]_sky130_fd_sc_hd__o221a_2_B2_B1_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[33]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a32o_2_X_A1  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a2bb2o_2_X_B2_sky130_fd_sc_hd__a22o_2_X_A1_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and4_2_X_B  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_hash_v_sky130_fd_sc_hd__a211o_2_X_A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_block_last_sky130_fd_sc_hd__a22o_2_B2_A1 (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout465_X (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[61]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[32]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[40]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[51]_sky130_fd_sc_hd__and3_2_A_B  (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_X (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_1_A  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_A  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout473_X (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[80]_sky130_fd_sc_hd__nand2_2_B_Y_sky130_fd_sc_hd__nor2_2_B_A_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__a31o_2_A3_A1  (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__or2_2_B_1_A  (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_B_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout476_X (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_B2_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nor2_2_A_1_B_sky130_fd_sc_hd__nand2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_B  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][0]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][9]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_q[1]_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout477_X (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_A  (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[3][13]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[10][30]_sky130_fd_sc_hd__and3_2_B_C_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[68]_sky130_fd_sc_hd__nor2_2_B_Y_sky130_fd_sc_hd__o22a_2_B1_A1_sky130_fd_sc_hd__nand2_2_Y_B  (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[25]_sky130_fd_sc_hd__a22o_2_X_A2_sky130_fd_sc_hd__and3_2_X_A  (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_c_buf[23]_sky130_fd_sc_hd__o311a_2_X_A1  (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[8][20]_sky130_fd_sc_hd__mux4_2_A0_S0  (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout476_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_X (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[201]_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.res_cnt_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__nor2_2_Y_A_sky130_fd_sc_hd__inv_2_Y_A  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.res_cnt_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_A  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o21a_2_X_A2_sky130_fd_sc_hd__a32o_2_X_B2  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.fsm_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__a221o_2_X_B2  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_hash_v_sky130_fd_sc_hd__a211o_2_X_C1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.shift_hash_q_sky130_fd_sc_hd__a21oi_2_A1_A2  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout480_X (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[207]_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[205]_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[175]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[141]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[171]_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C_B  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__a31o_2_A3_A2  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout484_X (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[104]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[112]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[57]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[97]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[65]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[34]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[42]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[50]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[82]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout483_A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout485_X (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[217]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[145]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[209]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[122]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.nn_q[0]_sky130_fd_sc_hd__nand2_2_A_B  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_block_first_sky130_fd_sc_hd__a22o_2_B2_A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[4]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[193]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[3]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[185]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout486_X (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[249]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[129]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[137]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout485_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[72]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[32]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[25]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout484_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout487_X (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[176]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[146]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__nor2_2_A_B  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[234]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[218]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[162]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[178]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[250]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__o32a_2_A2_A1  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout489_X (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout487_A (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout488_A (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[24]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[56]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[120]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[76]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[108]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[4]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout492_X (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[188]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[252]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[220]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[140]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[228]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[238]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[174]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[134]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout494_X (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout493_A (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[93]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[101]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[29]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[69]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout490_A (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout497_X (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[127]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout496_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[86]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[110]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout495_A (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout499_X (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[204]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[253]_sky130_fd_sc_hd__inv_2_A_Y_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[245]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[133]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout498_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[3]_sky130_fd_sc_hd__mux2_1_A1_S  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[246]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[254]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[158]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout500_X (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout499_A (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[125]_sky130_fd_sc_hd__nor2_2_B_A  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_hash[6]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[14]_sky130_fd_sc_hd__or2_2_B_A  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout497_A (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout509_X (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout508_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout504_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout502_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[48]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout505_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout520_X (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[203]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[235]_sky130_fd_sc_hd__and3_2_C_X_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[139]_sky130_fd_sc_hd__a31o_2_A3_B1  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[131]_sky130_fd_sc_hd__a22o_2_A1_B2_sky130_fd_sc_hd__nand2_2_Y_A  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[152]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[160]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[248]_sky130_fd_sc_hd__a22o_2_A1_B2  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[216]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[224]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[150]_sky130_fd_sc_hd__mux2_1_A0_S  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout524_X (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout520_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout523_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout522_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout519_A (.DIODE(net524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_X (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout532_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout537_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout526_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout530_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout539_X (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout524_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout509_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout516_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout511_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_X (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout599_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout590_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout561_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout546_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout550_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout579_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout614_X (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[41]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[42]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[49]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[50]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout613_A (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[56]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[4]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout615_X (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout614_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.cmd[5]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__and2_2_X_A  (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.kk_q[0]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__nor3_2_Y_B_sky130_fd_sc_hd__nand2_2_B_A  (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_X (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout618_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[60]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_io.m_config.ll_q[61]_sky130_fd_sc_hd__dfxtp_2_Q_D_sky130_fd_sc_hd__o211a_2_X_C1  (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout617_A (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload14_A (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[13][8]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][16]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[3][24]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[7][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[7][2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[8][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[3][16]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[8][18]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[8][26]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[15][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[15][2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[14][26]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[1][26]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[2][2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[6][26]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[2][18]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[2][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[1][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[0][2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[5][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_matrix[5][2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_X (.DIODE(clknet_leaf_17_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload29_A (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[14][8]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[136]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][0]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][0]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][0]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[18]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[128]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[19]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[130]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[0]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[1]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.g_idx_next[2]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[1]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][10]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[17]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_X (.DIODE(clknet_leaf_29_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[24]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[26]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.a_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[27]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][8]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][8]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[200]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[12][16]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][16]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[7][16]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[144]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][16]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[6][16]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[12]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[3]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[14]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.b_q[13]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][6]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.m_g.d_q[28]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[142]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[4][14]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.h_flat[206]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_m_blake2.m_hash256.v_q[5][6]_sky130_fd_sc_hd__dfxtp_2_Q_CLK  (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_X (.DIODE(clknet_leaf_48_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_A (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_clk_X (.DIODE(clknet_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_clk_A (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_clk_X (.DIODE(clknet_3_0_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_clk_A (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_clk_X (.DIODE(clknet_3_1_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_clk_A (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_clk_X (.DIODE(clknet_3_2_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload1_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_clk_A (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_clk_X (.DIODE(clknet_3_3_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload2_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_clk_A (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_clk_X (.DIODE(clknet_3_4_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload3_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_clk_A (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_clk_X (.DIODE(clknet_3_5_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload4_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_clk_A (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_clk_X (.DIODE(clknet_3_6_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload5_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_clk_A (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_clk_X (.DIODE(clknet_3_7_0_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\m_blake2.m_hash256.g_b[22]_sky130_fd_sc_hd__or2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__nand2_2_Y_A ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\m_blake2.m_hash256.g_b[9]_sky130_fd_sc_hd__and2_2_A_B_sky130_fd_sc_hd__xnor2_2_Y_A_sky130_fd_sc_hd__a21oi_2_Y_B1 ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\m_blake2.m_hash256.g_d[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\m_blake2.m_hash256.h_flat[56] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\m_blake2.m_hash256.m_g.a0[12]_sky130_fd_sc_hd__xor2_2_X_B_sky130_fd_sc_hd__or2_2_X_B ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\m_blake2.m_hash256.m_g.c_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\m_blake2.m_hash256.m_g.c_q[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\m_blake2.m_hash256.round_q[8]_sky130_fd_sc_hd__or4_2_A_X_sky130_fd_sc_hd__o31a_2_A3_X_sky130_fd_sc_hd__nand2b_2_A_N_Y_sky130_fd_sc_hd__nor2_2_B_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\m_blake2.m_hash256.v_q[9][5]_sky130_fd_sc_hd__and3_2_A_C_sky130_fd_sc_hd__nor2_2_B_1_Y ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\m_blake2.m_hash256.block_idx_plus_one_q[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\m_blake2.m_hash256.g_d[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\m_blake2.m_hash256.g_d[7] ));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_968 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1108 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1203 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1211 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1238 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1280 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1341 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1403 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1415 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1439 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1451 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1243 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1291 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1154 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1193 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1210 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1376 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_974 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1115 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1140 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1294 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1306 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1338 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1386 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1427 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1431 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1439 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1443 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1090 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1164 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1230 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1248 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1340 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1028 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1037 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1128 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1164 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1174 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1232 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1244 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1362 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1366 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1038 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1159 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1193 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1231 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1300 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1438 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1450 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1172 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1335 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1390 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1402 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1410 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1446 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1458 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1067 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1316 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1328 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1360 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1433 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1080 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1169 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1246 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1256 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1282 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1285 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1290 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1375 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1406 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1153 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1158 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1204 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1292 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1418 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1164 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1286 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1389 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1449 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1124 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1297 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1340 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1376 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1405 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1174 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1202 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_876 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1082 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1175 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1186 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1194 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1419 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1423 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_1447 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_1201 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1306 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1317 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1387 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1438 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1442 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1461 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1026 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1194 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1306 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1338 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1365 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1388 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1422 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1020 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1169 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1195 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1199 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1294 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1337 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1384 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1396 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1427 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1011 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1237 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1246 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1308 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1322 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1455 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_832 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1008 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1171 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1202 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1299 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1346 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1395 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1403 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1412 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1436 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1440 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1448 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1460 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1193 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1197 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1202 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1378 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1417 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1115 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_1123 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1168 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1190 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1358 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1370 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1394 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1258 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1291 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1340 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1345 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1357 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1403 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1435 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_1466 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1106 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1127 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1325 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1337 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1355 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1463 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1150 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1185 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1231 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1257 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1324 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1330 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1418 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_902 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1030 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1156 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1168 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1172 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1192 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1195 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1240 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1334 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1384 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1407 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1415 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1426 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_1434 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1467 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1154 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1199 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1246 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1280 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1361 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1408 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1432 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_862 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1023 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1155 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1173 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1315 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1337 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1347 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1423 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1427 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1133 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1174 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1240 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1276 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1289 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1364 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1376 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1398 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1421 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1434 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_611 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1114 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1205 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1259 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1272 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1279 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1325 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1382 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1427 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1429 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1438 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1134 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1268 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1274 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_973 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1158 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1170 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1174 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1330 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1388 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1402 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1414 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1418 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1466 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_988 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1031 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1043 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1208 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1220 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1228 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1356 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1419 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1465 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_616 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_952 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1002 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1039 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1181 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1334 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1349 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1393 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1420 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1427 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1467 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1047 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1081 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1173 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1185 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1208 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1312 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1396 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1455 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1172 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1259 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1307 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1346 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1390 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1429 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1042 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1156 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1179 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1409 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1433 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1443 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1452 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1466 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_494 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1015 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1142 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1176 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1214 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1265 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1360 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1438 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1464 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_935 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_972 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1118 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1190 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1214 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1278 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1317 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1436 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1100 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1108 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1163 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1192 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1217 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1254 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1272 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1313 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1404 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1448 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1460 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1468 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_798 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1124 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1208 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1218 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1263 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1327 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1352 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1375 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1399 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1401 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1066 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1214 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1234 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1315 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1321 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1385 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1463 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1116 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1135 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1204 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1226 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1286 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1358 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1366 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1410 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1454 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1468 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_844 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1176 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1250 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1257 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1313 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1319 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1400 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1412 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1427 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_1439 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1468 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_966 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1293 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1296 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1347 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1395 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1410 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1418 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_896 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1010 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1111 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1161 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1173 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1214 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1294 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_1313 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1335 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1467 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1123 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1204 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1318 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1330 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1399 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1420 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1444 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_956 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1084 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1147 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1165 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1203 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1275 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1456 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1266 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_1333 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1345 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1372 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1399 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1411 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1419 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1428 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1008 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1081 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1140 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1212 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1238 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1259 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1326 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1332 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1368 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1461 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_1326 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1334 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1359 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1377 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1218 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1256 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1270 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1290 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1315 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1338 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1346 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1355 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1371 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1416 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1427 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_1466 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1208 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1227 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1233 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1249 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1328 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1385 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1396 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1428 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1186 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1238 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1284 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1296 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1317 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1329 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1377 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1389 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1414 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1420 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1438 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1444 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_1454 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1462 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1468 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1146 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1200 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1208 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1230 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1237 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1325 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1361 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1408 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1427 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1442 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1182 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1229 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1279 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1358 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1397 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1411 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1437 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1459 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1467 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1293 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1349 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1438 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1466 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1034 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1173 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1306 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1341 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1366 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1398 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1468 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1074 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1153 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1184 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1224 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1283 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1289 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1351 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1399 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1452 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1467 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1105 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1113 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1180 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1228 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1234 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1297 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1315 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1335 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1371 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1405 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1456 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1468 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_906 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1173 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1185 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1230 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1233 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1241 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1254 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1269 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1297 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1327 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1386 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1405 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1065 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1181 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1225 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1237 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1258 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1289 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1338 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1342 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1382 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1424 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1458 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_1466 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1038 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1144 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1159 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1177 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1189 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1197 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1229 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1309 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1369 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1381 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1403 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1415 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1430 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1466 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_956 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1109 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1124 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1198 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1205 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1228 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1236 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1282 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1349 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1381 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1409 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1464 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1030 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1177 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1206 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1228 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1233 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1245 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1343 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1379 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1390 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1394 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1425 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1457 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_1466 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1068 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1239 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1336 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1378 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1382 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1402 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1427 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_1436 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1461 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1037 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1173 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1177 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1241 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1247 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1293 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1343 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_1352 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1360 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1399 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1424 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1438 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_1453 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_831 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_848 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1110 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1158 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1222 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1235 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1247 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1294 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1364 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_1454 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1464 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_415 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1039 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1163 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1213 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1218 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1235 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1248 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1265 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1286 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1295 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1325 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1349 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1426 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1465 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_952 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1221 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1277 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1296 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1300 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1305 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1312 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1333 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1341 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1365 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1401 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1426 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_990 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1166 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1188 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1246 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1287 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1371 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1397 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1409 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_1420 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1428 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1465 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_917 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1203 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1207 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1252 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1255 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1314 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1317 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1366 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1373 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1425 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1436 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1444 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1464 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1092 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1100 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1242 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1254 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1343 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1363 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1381 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1398 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1406 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1410 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1435 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1448 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1457 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1467 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_972 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1004 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1172 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1190 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1237 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1256 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1285 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1322 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1417 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1468 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1201 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1210 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1216 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1226 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1233 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1240 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1302 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1308 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1342 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1370 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1380 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1390 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1418 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1426 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1454 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1457 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1463 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1107 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1182 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1202 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1252 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1306 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1328 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1340 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1368 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1379 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1387 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1402 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1425 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_1466 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1112 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1262 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1333 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_1341 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1423 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1457 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1074 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1167 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1175 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1193 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1232 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1258 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1287 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1342 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1426 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1429 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1437 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1455 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1467 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1023 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1170 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1177 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1194 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1231 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1235 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1284 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1343 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1345 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1384 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1390 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1430 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1442 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1452 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1465 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1053 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1117 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1177 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1189 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1198 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1259 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1305 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1331 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1343 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1363 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1373 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1422 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1457 ();
 assign uio_oe[0] = net627;
 assign uio_oe[1] = net626;
 assign uio_oe[2] = net625;
 assign uio_oe[3] = net635;
 assign uio_oe[4] = net624;
 assign uio_oe[5] = net623;
 assign uio_oe[6] = net622;
 assign uio_oe[7] = net634;
 assign uio_out[0] = net633;
 assign uio_out[1] = net632;
 assign uio_out[2] = net631;
 assign uio_out[4] = net630;
 assign uio_out[5] = net629;
 assign uio_out[6] = net628;
endmodule
